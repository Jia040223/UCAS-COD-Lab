// ALU_AND
`STIMULI(3'd0, 32'hffffffff, 32'hffffffff)
`STIMULI(3'd0, 32'hfffffffe, 32'hffffffff)
`STIMULI(3'd0, 32'h80000001, 32'hffffffff)
`STIMULI(3'd0, 32'h80000000, 32'hffffffff)
`STIMULI(3'd0, 32'h7fffffff, 32'hffffffff)
`STIMULI(3'd0, 32'h00000002, 32'hffffffff)
`STIMULI(3'd0, 32'h00000001, 32'hffffffff)
`STIMULI(3'd0, 32'h00000000, 32'hffffffff)
`STIMULI(3'd0, 32'hffffffff, 32'hfffffffe)
`STIMULI(3'd0, 32'hfffffffe, 32'hfffffffe)
`STIMULI(3'd0, 32'h80000001, 32'hfffffffe)
`STIMULI(3'd0, 32'h80000000, 32'hfffffffe)
`STIMULI(3'd0, 32'h7fffffff, 32'hfffffffe)
`STIMULI(3'd0, 32'h00000002, 32'hfffffffe)
`STIMULI(3'd0, 32'h00000001, 32'hfffffffe)
`STIMULI(3'd0, 32'h00000000, 32'hfffffffe)
`STIMULI(3'd0, 32'hffffffff, 32'h80000001)
`STIMULI(3'd0, 32'hfffffffe, 32'h80000001)
`STIMULI(3'd0, 32'h80000001, 32'h80000001)
`STIMULI(3'd0, 32'h80000000, 32'h80000001)
`STIMULI(3'd0, 32'h7fffffff, 32'h80000001)
`STIMULI(3'd0, 32'h00000002, 32'h80000001)
`STIMULI(3'd0, 32'h00000001, 32'h80000001)
`STIMULI(3'd0, 32'h00000000, 32'h80000001)
`STIMULI(3'd0, 32'hffffffff, 32'h80000000)
`STIMULI(3'd0, 32'hfffffffe, 32'h80000000)
`STIMULI(3'd0, 32'h80000001, 32'h80000000)
`STIMULI(3'd0, 32'h80000000, 32'h80000000)
`STIMULI(3'd0, 32'h7fffffff, 32'h80000000)
`STIMULI(3'd0, 32'h00000002, 32'h80000000)
`STIMULI(3'd0, 32'h00000001, 32'h80000000)
`STIMULI(3'd0, 32'h00000000, 32'h80000000)
`STIMULI(3'd0, 32'hffffffff, 32'h7fffffff)
`STIMULI(3'd0, 32'hfffffffe, 32'h7fffffff)
`STIMULI(3'd0, 32'h80000001, 32'h7fffffff)
`STIMULI(3'd0, 32'h80000000, 32'h7fffffff)
`STIMULI(3'd0, 32'h7fffffff, 32'h7fffffff)
`STIMULI(3'd0, 32'h00000002, 32'h7fffffff)
`STIMULI(3'd0, 32'h00000001, 32'h7fffffff)
`STIMULI(3'd0, 32'h00000000, 32'h7fffffff)
`STIMULI(3'd0, 32'hffffffff, 32'h00000002)
`STIMULI(3'd0, 32'hfffffffe, 32'h00000002)
`STIMULI(3'd0, 32'h80000001, 32'h00000002)
`STIMULI(3'd0, 32'h80000000, 32'h00000002)
`STIMULI(3'd0, 32'h7fffffff, 32'h00000002)
`STIMULI(3'd0, 32'h00000002, 32'h00000002)
`STIMULI(3'd0, 32'h00000001, 32'h00000002)
`STIMULI(3'd0, 32'h00000000, 32'h00000002)
`STIMULI(3'd0, 32'hffffffff, 32'h00000001)
`STIMULI(3'd0, 32'hfffffffe, 32'h00000001)
`STIMULI(3'd0, 32'h80000001, 32'h00000001)
`STIMULI(3'd0, 32'h80000000, 32'h00000001)
`STIMULI(3'd0, 32'h7fffffff, 32'h00000001)
`STIMULI(3'd0, 32'h00000002, 32'h00000001)
`STIMULI(3'd0, 32'h00000001, 32'h00000001)
`STIMULI(3'd0, 32'h00000000, 32'h00000001)
`STIMULI(3'd0, 32'hffffffff, 32'h00000000)
`STIMULI(3'd0, 32'hfffffffe, 32'h00000000)
`STIMULI(3'd0, 32'h80000001, 32'h00000000)
`STIMULI(3'd0, 32'h80000000, 32'h00000000)
`STIMULI(3'd0, 32'h7fffffff, 32'h00000000)
`STIMULI(3'd0, 32'h00000002, 32'h00000000)
`STIMULI(3'd0, 32'h00000001, 32'h00000000)
`STIMULI(3'd0, 32'h00000000, 32'h00000000)
`STIMULI(3'd0, 32'h4b20e646, 32'h4da33da8)
`STIMULI(3'd0, 32'h5ab1862e, 32'hb8f81dca)
`STIMULI(3'd0, 32'h02b5a75c, 32'h7718eab3)
`STIMULI(3'd0, 32'h2c37a65a, 32'h4dd68da3)
`STIMULI(3'd0, 32'h44bc285c, 32'h86e92c89)
`STIMULI(3'd0, 32'h86ceab6d, 32'h4771cfb8)
`STIMULI(3'd0, 32'h7e02173c, 32'h330651c7)
`STIMULI(3'd0, 32'h15485d5b, 32'h42be3f98)
`STIMULI(3'd0, 32'h39ef7e50, 32'h1c1708c8)
`STIMULI(3'd0, 32'h8a300f51, 32'hb7f1958d)
`STIMULI(3'd0, 32'h4f1d5a90, 32'h1f786cac)
`STIMULI(3'd0, 32'h7aafd525, 32'h090cd8e0)
`STIMULI(3'd0, 32'hbb8f7575, 32'h04dfe476)
`STIMULI(3'd0, 32'h40fe6e6d, 32'h8aacd005)
`STIMULI(3'd0, 32'ha4585123, 32'hbbae4393)
`STIMULI(3'd0, 32'h13b9a8e5, 32'h5fe7c698)
`STIMULI(3'd0, 32'h408e2809, 32'h54b81753)
`STIMULI(3'd0, 32'h6a94969d, 32'h64e6792c)
`STIMULI(3'd0, 32'h90665ae6, 32'h7e4e3f82)
`STIMULI(3'd0, 32'h44ce3fc4, 32'h50f482ef)
`STIMULI(3'd0, 32'h530656d5, 32'h2f62d661)
`STIMULI(3'd0, 32'hb5dafc1c, 32'h636cb1bb)
`STIMULI(3'd0, 32'hadb115e4, 32'h7aa93be0)
`STIMULI(3'd0, 32'hb46134ab, 32'h00b76cb9)
`STIMULI(3'd0, 32'haa0c1242, 32'h6a3c30c7)
`STIMULI(3'd0, 32'h64241e75, 32'h57bd2826)
`STIMULI(3'd0, 32'h64e56ca7, 32'h98855320)
`STIMULI(3'd0, 32'h587494df, 32'h0ef17ee9)
`STIMULI(3'd0, 32'h82c183e7, 32'h3c98b354)
`STIMULI(3'd0, 32'h66aea70f, 32'h67a6f08e)
`STIMULI(3'd0, 32'h551e0674, 32'hbf233bef)
`STIMULI(3'd0, 32'h76986f78, 32'h57df8a5b)
`STIMULI(3'd0, 32'h7bbbef43, 32'h5d471687)
`STIMULI(3'd0, 32'hbf867aea, 32'h50d9f5b8)
`STIMULI(3'd0, 32'h1c6a5276, 32'hb61eea62)
`STIMULI(3'd0, 32'h28b98013, 32'h982641ba)
`STIMULI(3'd0, 32'h136600e9, 32'h683ffafd)
`STIMULI(3'd0, 32'h69003772, 32'hafd05360)
`STIMULI(3'd0, 32'h1e5ee55f, 32'h11b9b785)
`STIMULI(3'd0, 32'h47f6951a, 32'hb1c4e649)
`STIMULI(3'd0, 32'h79f9b283, 32'hb0f6cc8c)
`STIMULI(3'd0, 32'h619539a9, 32'h185897e2)
`STIMULI(3'd0, 32'h42b08411, 32'ha98bcec3)
`STIMULI(3'd0, 32'h4a1d7e2b, 32'h3caa3694)
`STIMULI(3'd0, 32'h5a829b4f, 32'h2bb2b7d4)
`STIMULI(3'd0, 32'h5502ce77, 32'h1d331f60)
`STIMULI(3'd0, 32'h553e8697, 32'h1f204ca2)
`STIMULI(3'd0, 32'h59dd55f5, 32'h2fc121e6)
`STIMULI(3'd0, 32'h4ad30477, 32'haee0246c)
`STIMULI(3'd0, 32'h4cf44147, 32'h20118b0e)
`STIMULI(3'd0, 32'h4e00710e, 32'ha6d1973c)
`STIMULI(3'd0, 32'h4fd2acf5, 32'h18d37585)
`STIMULI(3'd0, 32'h55b1bba8, 32'h9cc6ee3c)
`STIMULI(3'd0, 32'hb8e50094, 32'h23b22cb6)
`STIMULI(3'd0, 32'h43988578, 32'h88b7ad89)
`STIMULI(3'd0, 32'hbc85a23c, 32'h994a4120)
`STIMULI(3'd0, 32'ha57e9bc5, 32'h756aa2d0)
`STIMULI(3'd0, 32'h3cfc6dd6, 32'h6917213d)
`STIMULI(3'd0, 32'h7e225059, 32'h79821012)
`STIMULI(3'd0, 32'h8261625d, 32'ha3a0ec1e)
`STIMULI(3'd0, 32'h6eecb2e2, 32'h3f5dd033)
`STIMULI(3'd0, 32'h8cb80d5b, 32'h6d0f033b)
`STIMULI(3'd0, 32'hb8dfe046, 32'h8f196fb8)
`STIMULI(3'd0, 32'h10afef59, 32'h27cc9328)
`STIMULI(3'd0, 32'h4e773feb, 32'h1d67fcb4)
`STIMULI(3'd0, 32'h94db9664, 32'h07572031)
`STIMULI(3'd0, 32'h2c816c6c, 32'h258b85bd)
`STIMULI(3'd0, 32'haf23b35a, 32'h7af8ac58)
`STIMULI(3'd0, 32'h42f38272, 32'h43ff49be)

// ALU_OR
`STIMULI(3'd1, 32'hffffffff, 32'hffffffff)
`STIMULI(3'd1, 32'hfffffffe, 32'hffffffff)
`STIMULI(3'd1, 32'h80000001, 32'hffffffff)
`STIMULI(3'd1, 32'h80000000, 32'hffffffff)
`STIMULI(3'd1, 32'h7fffffff, 32'hffffffff)
`STIMULI(3'd1, 32'h00000002, 32'hffffffff)
`STIMULI(3'd1, 32'h00000001, 32'hffffffff)
`STIMULI(3'd1, 32'h00000000, 32'hffffffff)
`STIMULI(3'd1, 32'hffffffff, 32'hfffffffe)
`STIMULI(3'd1, 32'hfffffffe, 32'hfffffffe)
`STIMULI(3'd1, 32'h80000001, 32'hfffffffe)
`STIMULI(3'd1, 32'h80000000, 32'hfffffffe)
`STIMULI(3'd1, 32'h7fffffff, 32'hfffffffe)
`STIMULI(3'd1, 32'h00000002, 32'hfffffffe)
`STIMULI(3'd1, 32'h00000001, 32'hfffffffe)
`STIMULI(3'd1, 32'h00000000, 32'hfffffffe)
`STIMULI(3'd1, 32'hffffffff, 32'h80000001)
`STIMULI(3'd1, 32'hfffffffe, 32'h80000001)
`STIMULI(3'd1, 32'h80000001, 32'h80000001)
`STIMULI(3'd1, 32'h80000000, 32'h80000001)
`STIMULI(3'd1, 32'h7fffffff, 32'h80000001)
`STIMULI(3'd1, 32'h00000002, 32'h80000001)
`STIMULI(3'd1, 32'h00000001, 32'h80000001)
`STIMULI(3'd1, 32'h00000000, 32'h80000001)
`STIMULI(3'd1, 32'hffffffff, 32'h80000000)
`STIMULI(3'd1, 32'hfffffffe, 32'h80000000)
`STIMULI(3'd1, 32'h80000001, 32'h80000000)
`STIMULI(3'd1, 32'h80000000, 32'h80000000)
`STIMULI(3'd1, 32'h7fffffff, 32'h80000000)
`STIMULI(3'd1, 32'h00000002, 32'h80000000)
`STIMULI(3'd1, 32'h00000001, 32'h80000000)
`STIMULI(3'd1, 32'h00000000, 32'h80000000)
`STIMULI(3'd1, 32'hffffffff, 32'h7fffffff)
`STIMULI(3'd1, 32'hfffffffe, 32'h7fffffff)
`STIMULI(3'd1, 32'h80000001, 32'h7fffffff)
`STIMULI(3'd1, 32'h80000000, 32'h7fffffff)
`STIMULI(3'd1, 32'h7fffffff, 32'h7fffffff)
`STIMULI(3'd1, 32'h00000002, 32'h7fffffff)
`STIMULI(3'd1, 32'h00000001, 32'h7fffffff)
`STIMULI(3'd1, 32'h00000000, 32'h7fffffff)
`STIMULI(3'd1, 32'hffffffff, 32'h00000002)
`STIMULI(3'd1, 32'hfffffffe, 32'h00000002)
`STIMULI(3'd1, 32'h80000001, 32'h00000002)
`STIMULI(3'd1, 32'h80000000, 32'h00000002)
`STIMULI(3'd1, 32'h7fffffff, 32'h00000002)
`STIMULI(3'd1, 32'h00000002, 32'h00000002)
`STIMULI(3'd1, 32'h00000001, 32'h00000002)
`STIMULI(3'd1, 32'h00000000, 32'h00000002)
`STIMULI(3'd1, 32'hffffffff, 32'h00000001)
`STIMULI(3'd1, 32'hfffffffe, 32'h00000001)
`STIMULI(3'd1, 32'h80000001, 32'h00000001)
`STIMULI(3'd1, 32'h80000000, 32'h00000001)
`STIMULI(3'd1, 32'h7fffffff, 32'h00000001)
`STIMULI(3'd1, 32'h00000002, 32'h00000001)
`STIMULI(3'd1, 32'h00000001, 32'h00000001)
`STIMULI(3'd1, 32'h00000000, 32'h00000001)
`STIMULI(3'd1, 32'hffffffff, 32'h00000000)
`STIMULI(3'd1, 32'hfffffffe, 32'h00000000)
`STIMULI(3'd1, 32'h80000001, 32'h00000000)
`STIMULI(3'd1, 32'h80000000, 32'h00000000)
`STIMULI(3'd1, 32'h7fffffff, 32'h00000000)
`STIMULI(3'd1, 32'h00000002, 32'h00000000)
`STIMULI(3'd1, 32'h00000001, 32'h00000000)
`STIMULI(3'd1, 32'h00000000, 32'h00000000)
`STIMULI(3'd1, 32'h024fcc89, 32'h6f74eede)
`STIMULI(3'd1, 32'h698acf7b, 32'h31737fe3)
`STIMULI(3'd1, 32'h6a6d9b36, 32'h2c7e51ed)
`STIMULI(3'd1, 32'h7572c9a1, 32'h6cbd67c0)
`STIMULI(3'd1, 32'h9bf340cc, 32'h5efd991d)
`STIMULI(3'd1, 32'h1e30e7a3, 32'h0660dc02)
`STIMULI(3'd1, 32'h0b7beb0a, 32'h93a3b145)
`STIMULI(3'd1, 32'h731e43c2, 32'h276f2bd6)
`STIMULI(3'd1, 32'h72a14a62, 32'h914f2b66)
`STIMULI(3'd1, 32'hadd007d9, 32'h7e1d356c)
`STIMULI(3'd1, 32'ha4f2dcab, 32'h20ee4b9b)
`STIMULI(3'd1, 32'ha58c6143, 32'h9794270d)
`STIMULI(3'd1, 32'h323d7701, 32'h535c691c)
`STIMULI(3'd1, 32'h15b15c79, 32'h573053ac)
`STIMULI(3'd1, 32'h744ab4b7, 32'h3b3dbdbc)
`STIMULI(3'd1, 32'h6ec47ab9, 32'ha6882bb9)
`STIMULI(3'd1, 32'h0e9a26d8, 32'h8475d733)
`STIMULI(3'd1, 32'h7db87f65, 32'h82e4db90)
`STIMULI(3'd1, 32'h3fb394ef, 32'h6c7cfa1f)
`STIMULI(3'd1, 32'ha96d0749, 32'h4e4dbbc8)
`STIMULI(3'd1, 32'h70f2d152, 32'h272586ae)
`STIMULI(3'd1, 32'h51329758, 32'h30a66641)
`STIMULI(3'd1, 32'h13a280cd, 32'h7a9f9ea1)
`STIMULI(3'd1, 32'h7ef42209, 32'h0495521f)
`STIMULI(3'd1, 32'h21c5254f, 32'h5026b961)
`STIMULI(3'd1, 32'hb53bb861, 32'hb567a61d)
`STIMULI(3'd1, 32'h4ac65802, 32'h342fda6a)
`STIMULI(3'd1, 32'h39fcf83c, 32'h6c8b7d52)
`STIMULI(3'd1, 32'h845693cc, 32'h6f38b09d)
`STIMULI(3'd1, 32'ha1f3236f, 32'h4f1cebce)
`STIMULI(3'd1, 32'ha3688b08, 32'h5bf01bab)
`STIMULI(3'd1, 32'h3ba86920, 32'ha7bf1ed4)
`STIMULI(3'd1, 32'h4b28cc49, 32'h5d9b8c8f)
`STIMULI(3'd1, 32'h76dc0aa2, 32'h6e915751)
`STIMULI(3'd1, 32'hb98ba83b, 32'hb28473c3)
`STIMULI(3'd1, 32'h96507625, 32'h84b47484)
`STIMULI(3'd1, 32'h10200052, 32'h0d2c80c7)
`STIMULI(3'd1, 32'h7345cbd5, 32'h49aba88d)
`STIMULI(3'd1, 32'h3fb0f48a, 32'h899641fa)
`STIMULI(3'd1, 32'h4e601d11, 32'h4fd0f4dd)
`STIMULI(3'd1, 32'h16c2c2c1, 32'h41a5e8e6)
`STIMULI(3'd1, 32'h197c9d6a, 32'h5673b74c)
`STIMULI(3'd1, 32'h4b3c2ae0, 32'h67dcba7c)
`STIMULI(3'd1, 32'ha644ac29, 32'h61feeda2)
`STIMULI(3'd1, 32'h2982a362, 32'h3fc14993)
`STIMULI(3'd1, 32'hb872a4ee, 32'h74bece43)
`STIMULI(3'd1, 32'h279e040f, 32'h5eb75117)
`STIMULI(3'd1, 32'h56bdbbe5, 32'h5120a772)
`STIMULI(3'd1, 32'h1e789aaa, 32'h8f3060d3)
`STIMULI(3'd1, 32'h45df75b5, 32'h46169eba)
`STIMULI(3'd1, 32'h6de7b1ea, 32'h9c9d319a)
`STIMULI(3'd1, 32'h9737462c, 32'h0c604c94)
`STIMULI(3'd1, 32'habcd926d, 32'h5d16bbe1)
`STIMULI(3'd1, 32'h5276eb4e, 32'h99b54457)
`STIMULI(3'd1, 32'h79b3ed7b, 32'h69ae317a)
`STIMULI(3'd1, 32'h261590eb, 32'ha5817fe8)
`STIMULI(3'd1, 32'h46c4ed5b, 32'h788c7c3a)
`STIMULI(3'd1, 32'hbf36c43f, 32'h4078dad6)
`STIMULI(3'd1, 32'h623aadb4, 32'h654c552a)
`STIMULI(3'd1, 32'h65fa5abe, 32'ha8ff9b10)
`STIMULI(3'd1, 32'h5dd8d164, 32'h25311efd)
`STIMULI(3'd1, 32'h697875e6, 32'h40137f19)
`STIMULI(3'd1, 32'h8a7d7428, 32'h4f72d0a5)
`STIMULI(3'd1, 32'h69131a29, 32'h6856458c)
`STIMULI(3'd1, 32'h74a3efa2, 32'h528b900f)
`STIMULI(3'd1, 32'h2869c4a5, 32'h7f2163ca)
`STIMULI(3'd1, 32'h21fe60b4, 32'h117cdece)
`STIMULI(3'd1, 32'h6777a957, 32'h96a25057)
`STIMULI(3'd1, 32'h64086ede, 32'h0fe16dfc)

// ALU_ADD
`STIMULI(3'd2, 32'hffffffff, 32'hffffffff)
`STIMULI(3'd2, 32'hfffffffe, 32'hffffffff)
`STIMULI(3'd2, 32'h80000001, 32'hffffffff)
`STIMULI(3'd2, 32'h80000000, 32'hffffffff)
`STIMULI(3'd2, 32'h7fffffff, 32'hffffffff)
`STIMULI(3'd2, 32'h00000002, 32'hffffffff)
`STIMULI(3'd2, 32'h00000001, 32'hffffffff)
`STIMULI(3'd2, 32'h00000000, 32'hffffffff)
`STIMULI(3'd2, 32'hffffffff, 32'hfffffffe)
`STIMULI(3'd2, 32'hfffffffe, 32'hfffffffe)
`STIMULI(3'd2, 32'h80000001, 32'hfffffffe)
`STIMULI(3'd2, 32'h80000000, 32'hfffffffe)
`STIMULI(3'd2, 32'h7fffffff, 32'hfffffffe)
`STIMULI(3'd2, 32'h00000002, 32'hfffffffe)
`STIMULI(3'd2, 32'h00000001, 32'hfffffffe)
`STIMULI(3'd2, 32'h00000000, 32'hfffffffe)
`STIMULI(3'd2, 32'hffffffff, 32'h80000001)
`STIMULI(3'd2, 32'hfffffffe, 32'h80000001)
`STIMULI(3'd2, 32'h80000001, 32'h80000001)
`STIMULI(3'd2, 32'h80000000, 32'h80000001)
`STIMULI(3'd2, 32'h7fffffff, 32'h80000001)
`STIMULI(3'd2, 32'h00000002, 32'h80000001)
`STIMULI(3'd2, 32'h00000001, 32'h80000001)
`STIMULI(3'd2, 32'h00000000, 32'h80000001)
`STIMULI(3'd2, 32'hffffffff, 32'h80000000)
`STIMULI(3'd2, 32'hfffffffe, 32'h80000000)
`STIMULI(3'd2, 32'h80000001, 32'h80000000)
`STIMULI(3'd2, 32'h80000000, 32'h80000000)
`STIMULI(3'd2, 32'h7fffffff, 32'h80000000)
`STIMULI(3'd2, 32'h00000002, 32'h80000000)
`STIMULI(3'd2, 32'h00000001, 32'h80000000)
`STIMULI(3'd2, 32'h00000000, 32'h80000000)
`STIMULI(3'd2, 32'hffffffff, 32'h7fffffff)
`STIMULI(3'd2, 32'hfffffffe, 32'h7fffffff)
`STIMULI(3'd2, 32'h80000001, 32'h7fffffff)
`STIMULI(3'd2, 32'h80000000, 32'h7fffffff)
`STIMULI(3'd2, 32'h7fffffff, 32'h7fffffff)
`STIMULI(3'd2, 32'h00000002, 32'h7fffffff)
`STIMULI(3'd2, 32'h00000001, 32'h7fffffff)
`STIMULI(3'd2, 32'h00000000, 32'h7fffffff)
`STIMULI(3'd2, 32'hffffffff, 32'h00000002)
`STIMULI(3'd2, 32'hfffffffe, 32'h00000002)
`STIMULI(3'd2, 32'h80000001, 32'h00000002)
`STIMULI(3'd2, 32'h80000000, 32'h00000002)
`STIMULI(3'd2, 32'h7fffffff, 32'h00000002)
`STIMULI(3'd2, 32'h00000002, 32'h00000002)
`STIMULI(3'd2, 32'h00000001, 32'h00000002)
`STIMULI(3'd2, 32'h00000000, 32'h00000002)
`STIMULI(3'd2, 32'hffffffff, 32'h00000001)
`STIMULI(3'd2, 32'hfffffffe, 32'h00000001)
`STIMULI(3'd2, 32'h80000001, 32'h00000001)
`STIMULI(3'd2, 32'h80000000, 32'h00000001)
`STIMULI(3'd2, 32'h7fffffff, 32'h00000001)
`STIMULI(3'd2, 32'h00000002, 32'h00000001)
`STIMULI(3'd2, 32'h00000001, 32'h00000001)
`STIMULI(3'd2, 32'h00000000, 32'h00000001)
`STIMULI(3'd2, 32'hffffffff, 32'h00000000)
`STIMULI(3'd2, 32'hfffffffe, 32'h00000000)
`STIMULI(3'd2, 32'h80000001, 32'h00000000)
`STIMULI(3'd2, 32'h80000000, 32'h00000000)
`STIMULI(3'd2, 32'h7fffffff, 32'h00000000)
`STIMULI(3'd2, 32'h00000002, 32'h00000000)
`STIMULI(3'd2, 32'h00000001, 32'h00000000)
`STIMULI(3'd2, 32'h00000000, 32'h00000000)
`STIMULI(3'd2, 32'h15c3b421, 32'h0606cf92)
`STIMULI(3'd2, 32'ha15e4ccb, 32'h7d3b5d78)
`STIMULI(3'd2, 32'h1ca91fe9, 32'h8566bba9)
`STIMULI(3'd2, 32'h8d1ccb75, 32'hb26cd40b)
`STIMULI(3'd2, 32'h0b6d8b3b, 32'hae7b1840)
`STIMULI(3'd2, 32'h2fa83183, 32'ha816ab25)
`STIMULI(3'd2, 32'hb3e1d3e9, 32'h3cc4fcf8)
`STIMULI(3'd2, 32'h5a837f30, 32'h3f4f5f24)
`STIMULI(3'd2, 32'h6b401538, 32'h0a2bb0b3)
`STIMULI(3'd2, 32'h67660a49, 32'h1f21e921)
`STIMULI(3'd2, 32'h46f0adac, 32'h41e98979)
`STIMULI(3'd2, 32'h5e714846, 32'h3230c2e4)
`STIMULI(3'd2, 32'h4c153a2d, 32'h45d7528f)
`STIMULI(3'd2, 32'h5152ac06, 32'h9305e7d9)
`STIMULI(3'd2, 32'h87c0dc09, 32'hafc3f44c)
`STIMULI(3'd2, 32'h4536aabd, 32'h53d61636)
`STIMULI(3'd2, 32'h759b46db, 32'h168956c3)
`STIMULI(3'd2, 32'h66dbfe0f, 32'h7d5c22e4)
`STIMULI(3'd2, 32'h464d4b0f, 32'h2c12a8cc)
`STIMULI(3'd2, 32'h5132391a, 32'hbbe891eb)
`STIMULI(3'd2, 32'h429bff90, 32'h380e3729)
`STIMULI(3'd2, 32'h3944b4cf, 32'h08e94a9f)
`STIMULI(3'd2, 32'h6420dff6, 32'h8a76edea)
`STIMULI(3'd2, 32'h44d1dc8a, 32'ha6bcdf86)
`STIMULI(3'd2, 32'h42852513, 32'h7e16915a)
`STIMULI(3'd2, 32'h2fa62a25, 32'h26a60509)
`STIMULI(3'd2, 32'h888d7f44, 32'h747806b0)
`STIMULI(3'd2, 32'h4d62e48f, 32'h4b12a457)
`STIMULI(3'd2, 32'h728e980a, 32'h7d090eb5)
`STIMULI(3'd2, 32'h71b8a961, 32'h7b1c174e)
`STIMULI(3'd2, 32'h71811565, 32'h3f1b8df0)
`STIMULI(3'd2, 32'h462ebba5, 32'h640fad6f)
`STIMULI(3'd2, 32'h3c249ca5, 32'h37e76506)
`STIMULI(3'd2, 32'h5f2bc4bd, 32'h2da5b20a)
`STIMULI(3'd2, 32'h7702f2f7, 32'h255a8062)
`STIMULI(3'd2, 32'h11b55f79, 32'h33278f9c)
`STIMULI(3'd2, 32'h5d41e569, 32'h70e12436)
`STIMULI(3'd2, 32'h60cd41a7, 32'h5444d860)
`STIMULI(3'd2, 32'h963ba499, 32'h7282a120)
`STIMULI(3'd2, 32'h076c67fc, 32'h737d8a02)
`STIMULI(3'd2, 32'h6363c557, 32'h6839a9a3)
`STIMULI(3'd2, 32'h47c26262, 32'h799f69f0)
`STIMULI(3'd2, 32'h5abc4ac4, 32'h4f2eca5e)
`STIMULI(3'd2, 32'h6d1cf3f2, 32'hbe20101b)
`STIMULI(3'd2, 32'hb7687402, 32'hb4df5654)
`STIMULI(3'd2, 32'hb7bf7a0b, 32'h9224bec6)
`STIMULI(3'd2, 32'h040e20b2, 32'ha4dc6dfd)
`STIMULI(3'd2, 32'h5044cee1, 32'h3b7694b4)
`STIMULI(3'd2, 32'h59bbc451, 32'h880448ec)
`STIMULI(3'd2, 32'h4d9b537a, 32'h5dc9e503)
`STIMULI(3'd2, 32'hace0b6e9, 32'h1de0225b)
`STIMULI(3'd2, 32'h994079b8, 32'h869c7b3a)
`STIMULI(3'd2, 32'h25e46b47, 32'h66dbcd32)
`STIMULI(3'd2, 32'h6466603d, 32'h52c52230)
`STIMULI(3'd2, 32'h84bbef8e, 32'h7da6d9f5)
`STIMULI(3'd2, 32'h59619d6a, 32'h2aa05ad5)
`STIMULI(3'd2, 32'h6482a728, 32'hbdc7fda8)
`STIMULI(3'd2, 32'h7d657d06, 32'h693e96b6)
`STIMULI(3'd2, 32'h3b6ed79d, 32'h56c71a70)
`STIMULI(3'd2, 32'h13def18b, 32'h1ff17ec5)
`STIMULI(3'd2, 32'h148f1818, 32'h11446e91)
`STIMULI(3'd2, 32'h0930157b, 32'h4ffdefb6)
`STIMULI(3'd2, 32'h680b8902, 32'h9d0f0707)
`STIMULI(3'd2, 32'h6fef6e7b, 32'h7c9aa11a)
`STIMULI(3'd2, 32'h2e537598, 32'h791f83f7)
`STIMULI(3'd2, 32'h4c9890d0, 32'h165efe9a)
`STIMULI(3'd2, 32'h962e8afe, 32'hbc87ff4c)
`STIMULI(3'd2, 32'h92f99fb5, 32'h44820096)
`STIMULI(3'd2, 32'hb5a78343, 32'h5f923085)

// ALU_SUB
`STIMULI(3'd6, 32'h5ae0ff31, 32'h4bd60e41)
`STIMULI(3'd6, 32'hffffffff, 32'hffffffff)
`STIMULI(3'd6, 32'hfffffffe, 32'hffffffff)
`STIMULI(3'd6, 32'h80000001, 32'hffffffff)
`STIMULI(3'd6, 32'h80000000, 32'hffffffff)
`STIMULI(3'd6, 32'h7fffffff, 32'hffffffff)
`STIMULI(3'd6, 32'h00000002, 32'hffffffff)
`STIMULI(3'd6, 32'h00000001, 32'hffffffff)
`STIMULI(3'd6, 32'h00000000, 32'hffffffff)
`STIMULI(3'd6, 32'hffffffff, 32'hfffffffe)
`STIMULI(3'd6, 32'hfffffffe, 32'hfffffffe)
`STIMULI(3'd6, 32'h80000001, 32'hfffffffe)
`STIMULI(3'd6, 32'h80000000, 32'hfffffffe)
`STIMULI(3'd6, 32'h7fffffff, 32'hfffffffe)
`STIMULI(3'd6, 32'h00000002, 32'hfffffffe)
`STIMULI(3'd6, 32'h00000001, 32'hfffffffe)
`STIMULI(3'd6, 32'h00000000, 32'hfffffffe)
`STIMULI(3'd6, 32'hffffffff, 32'h80000001)
`STIMULI(3'd6, 32'hfffffffe, 32'h80000001)
`STIMULI(3'd6, 32'h80000001, 32'h80000001)
`STIMULI(3'd6, 32'h80000000, 32'h80000001)
`STIMULI(3'd6, 32'h7fffffff, 32'h80000001)
`STIMULI(3'd6, 32'h00000002, 32'h80000001)
`STIMULI(3'd6, 32'h00000001, 32'h80000001)
`STIMULI(3'd6, 32'h00000000, 32'h80000001)
`STIMULI(3'd6, 32'hffffffff, 32'h80000000)
`STIMULI(3'd6, 32'hfffffffe, 32'h80000000)
`STIMULI(3'd6, 32'h80000001, 32'h80000000)
`STIMULI(3'd6, 32'h80000000, 32'h80000000)
`STIMULI(3'd6, 32'h7fffffff, 32'h80000000)
`STIMULI(3'd6, 32'h00000002, 32'h80000000)
`STIMULI(3'd6, 32'h00000001, 32'h80000000)
`STIMULI(3'd6, 32'h00000000, 32'h80000000)
`STIMULI(3'd6, 32'hffffffff, 32'h7fffffff)
`STIMULI(3'd6, 32'hfffffffe, 32'h7fffffff)
`STIMULI(3'd6, 32'h80000001, 32'h7fffffff)
`STIMULI(3'd6, 32'h80000000, 32'h7fffffff)
`STIMULI(3'd6, 32'h7fffffff, 32'h7fffffff)
`STIMULI(3'd6, 32'h00000002, 32'h7fffffff)
`STIMULI(3'd6, 32'h00000001, 32'h7fffffff)
`STIMULI(3'd6, 32'h00000000, 32'h7fffffff)
`STIMULI(3'd6, 32'hffffffff, 32'h00000002)
`STIMULI(3'd6, 32'hfffffffe, 32'h00000002)
`STIMULI(3'd6, 32'h80000001, 32'h00000002)
`STIMULI(3'd6, 32'h80000000, 32'h00000002)
`STIMULI(3'd6, 32'h7fffffff, 32'h00000002)
`STIMULI(3'd6, 32'h00000002, 32'h00000002)
`STIMULI(3'd6, 32'h00000001, 32'h00000002)
`STIMULI(3'd6, 32'h00000000, 32'h00000002)
`STIMULI(3'd6, 32'hffffffff, 32'h00000001)
`STIMULI(3'd6, 32'hfffffffe, 32'h00000001)
`STIMULI(3'd6, 32'h80000001, 32'h00000001)
`STIMULI(3'd6, 32'h80000000, 32'h00000001)
`STIMULI(3'd6, 32'h7fffffff, 32'h00000001)
`STIMULI(3'd6, 32'h00000002, 32'h00000001)
`STIMULI(3'd6, 32'h00000001, 32'h00000001)
`STIMULI(3'd6, 32'h00000000, 32'h00000001)
`STIMULI(3'd6, 32'hffffffff, 32'h00000000)
`STIMULI(3'd6, 32'hfffffffe, 32'h00000000)
`STIMULI(3'd6, 32'h80000001, 32'h00000000)
`STIMULI(3'd6, 32'h80000000, 32'h00000000)
`STIMULI(3'd6, 32'h7fffffff, 32'h00000000)
`STIMULI(3'd6, 32'h00000002, 32'h00000000)
`STIMULI(3'd6, 32'h00000001, 32'h00000000)
`STIMULI(3'd6, 32'h00000000, 32'h00000000)
`STIMULI(3'd6, 32'h1c1a2fd1, 32'h6dda9ee6)
`STIMULI(3'd6, 32'h10580ed7, 32'h51c1b314)
`STIMULI(3'd6, 32'h4d6ccf6b, 32'h6b390e08)
`STIMULI(3'd6, 32'h1d97c155, 32'h6986ff3d)
`STIMULI(3'd6, 32'h5913acee, 32'hadefd02d)
`STIMULI(3'd6, 32'h3b48b251, 32'ha6807c5a)
`STIMULI(3'd6, 32'h1928de35, 32'h58e073a7)
`STIMULI(3'd6, 32'h90077b97, 32'h723c8b24)
`STIMULI(3'd6, 32'h86d043d4, 32'h4b502de8)
`STIMULI(3'd6, 32'h98bd077e, 32'h1ff92209)
`STIMULI(3'd6, 32'h2430a18f, 32'ha8c48315)
`STIMULI(3'd6, 32'h1235ad2d, 32'h2b00e563)
`STIMULI(3'd6, 32'h7414b0fd, 32'h2af2b4ab)
`STIMULI(3'd6, 32'h4afa076d, 32'h9845528d)
`STIMULI(3'd6, 32'h53b737c0, 32'h5d2fb49a)
`STIMULI(3'd6, 32'h434637f0, 32'h47cbe8be)
`STIMULI(3'd6, 32'h88226946, 32'h0e403f5d)
`STIMULI(3'd6, 32'h60113b4b, 32'h5bd9a106)
`STIMULI(3'd6, 32'h6b6ff3f8, 32'h2357733b)
`STIMULI(3'd6, 32'h23a589c4, 32'h73925d3e)
`STIMULI(3'd6, 32'hb197b299, 32'h03b6c50f)
`STIMULI(3'd6, 32'h4f6bfe44, 32'h9d07a691)
`STIMULI(3'd6, 32'ha70e384b, 32'h73118809)
`STIMULI(3'd6, 32'h909a03cf, 32'h58a5eae4)
`STIMULI(3'd6, 32'h76c84d18, 32'h60060213)
`STIMULI(3'd6, 32'h75ad9175, 32'h1dd68563)
`STIMULI(3'd6, 32'h53178a1c, 32'h86479544)
`STIMULI(3'd6, 32'h767c7047, 32'h49dfd735)
`STIMULI(3'd6, 32'h664d9757, 32'h6c2a01bc)
`STIMULI(3'd6, 32'h67b65c98, 32'hb9652174)
`STIMULI(3'd6, 32'h72719700, 32'h5e32cce0)
`STIMULI(3'd6, 32'h8344f8a9, 32'h58bf2e58)
`STIMULI(3'd6, 32'h4a5cce9c, 32'h6afb5541)
`STIMULI(3'd6, 32'h92244fcc, 32'hbcce659d)
`STIMULI(3'd6, 32'h492e2221, 32'h95694875)
`STIMULI(3'd6, 32'h958d93f5, 32'h938af0be)
`STIMULI(3'd6, 32'h00649db6, 32'ha7b1e3c1)
`STIMULI(3'd6, 32'h5059565b, 32'h4992bfd8)
`STIMULI(3'd6, 32'hbd1b2c36, 32'h65e6ea50)
`STIMULI(3'd6, 32'h5d1db096, 32'h3d7fc9ec)
`STIMULI(3'd6, 32'h8d98ce11, 32'had7706f1)
`STIMULI(3'd6, 32'h071289c4, 32'h4ab3fa47)
`STIMULI(3'd6, 32'h935df141, 32'h64303a5a)
`STIMULI(3'd6, 32'h0833c433, 32'ha0f6bf52)
`STIMULI(3'd6, 32'h11a7414b, 32'h8f464df8)
`STIMULI(3'd6, 32'h6baab999, 32'h2505328c)
`STIMULI(3'd6, 32'h73768852, 32'h73de7dcc)
`STIMULI(3'd6, 32'h45fbf1de, 32'h851dc99e)
`STIMULI(3'd6, 32'h0324cbc4, 32'h31a6ab77)
`STIMULI(3'd6, 32'h2a22fc2a, 32'h769b5417)
`STIMULI(3'd6, 32'ha5852944, 32'h701eee09)
`STIMULI(3'd6, 32'h7bb91db5, 32'h28a9f508)
`STIMULI(3'd6, 32'h21c59980, 32'h25dc19df)
`STIMULI(3'd6, 32'h1f45491f, 32'h474ac2c4)
`STIMULI(3'd6, 32'h15fb07e8, 32'h1afe66d4)
`STIMULI(3'd6, 32'h6ff4b7cd, 32'hb7c0a169)
`STIMULI(3'd6, 32'h40da80b4, 32'h0f3a00ec)
`STIMULI(3'd6, 32'h7f0b642d, 32'h56d5889c)
`STIMULI(3'd6, 32'haa3867c1, 32'h6f001bfa)
`STIMULI(3'd6, 32'h0e962a05, 32'h6b12e875)
`STIMULI(3'd6, 32'h7e3a1ce7, 32'h8da18e33)
`STIMULI(3'd6, 32'h41e87111, 32'ha87284a8)
`STIMULI(3'd6, 32'h7ca1aa2d, 32'h507e9b17)
`STIMULI(3'd6, 32'h93856d1d, 32'h7adbc714)
`STIMULI(3'd6, 32'h5e20294a, 32'h556dde2e)
`STIMULI(3'd6, 32'h234e4bbc, 32'h5ac1d377)
`STIMULI(3'd6, 32'h25ec7945, 32'h36d3b8d9)
`STIMULI(3'd6, 32'h559d9a8c, 32'h040ca28f)
`STIMULI(3'd6, 32'h8c419708, 32'h78ebe648)

// ALU_SLT
`STIMULI(3'd7, 32'hffffffff, 32'hffffffff)
`STIMULI(3'd7, 32'hfffffffe, 32'hffffffff)
`STIMULI(3'd7, 32'h80000001, 32'hffffffff)
`STIMULI(3'd7, 32'h80000000, 32'hffffffff)
`STIMULI(3'd7, 32'h7fffffff, 32'hffffffff)
`STIMULI(3'd7, 32'h00000002, 32'hffffffff)
`STIMULI(3'd7, 32'h00000001, 32'hffffffff)
`STIMULI(3'd7, 32'h00000000, 32'hffffffff)
`STIMULI(3'd7, 32'hffffffff, 32'hfffffffe)
`STIMULI(3'd7, 32'hfffffffe, 32'hfffffffe)
`STIMULI(3'd7, 32'h80000001, 32'hfffffffe)
`STIMULI(3'd7, 32'h80000000, 32'hfffffffe)
`STIMULI(3'd7, 32'h7fffffff, 32'hfffffffe)
`STIMULI(3'd7, 32'h00000002, 32'hfffffffe)
`STIMULI(3'd7, 32'h00000001, 32'hfffffffe)
`STIMULI(3'd7, 32'h00000000, 32'hfffffffe)
`STIMULI(3'd7, 32'hffffffff, 32'h80000001)
`STIMULI(3'd7, 32'hfffffffe, 32'h80000001)
`STIMULI(3'd7, 32'h80000001, 32'h80000001)
`STIMULI(3'd7, 32'h80000000, 32'h80000001)
`STIMULI(3'd7, 32'h7fffffff, 32'h80000001)
`STIMULI(3'd7, 32'h00000002, 32'h80000001)
`STIMULI(3'd7, 32'h00000001, 32'h80000001)
`STIMULI(3'd7, 32'h00000000, 32'h80000001)
`STIMULI(3'd7, 32'hffffffff, 32'h80000000)
`STIMULI(3'd7, 32'hfffffffe, 32'h80000000)
`STIMULI(3'd7, 32'h80000001, 32'h80000000)
`STIMULI(3'd7, 32'h80000000, 32'h80000000)
`STIMULI(3'd7, 32'h7fffffff, 32'h80000000)
`STIMULI(3'd7, 32'h00000002, 32'h80000000)
`STIMULI(3'd7, 32'h00000001, 32'h80000000)
`STIMULI(3'd7, 32'h00000000, 32'h80000000)
`STIMULI(3'd7, 32'hffffffff, 32'h7fffffff)
`STIMULI(3'd7, 32'hfffffffe, 32'h7fffffff)
`STIMULI(3'd7, 32'h80000001, 32'h7fffffff)
`STIMULI(3'd7, 32'h80000000, 32'h7fffffff)
`STIMULI(3'd7, 32'h7fffffff, 32'h7fffffff)
`STIMULI(3'd7, 32'h00000002, 32'h7fffffff)
`STIMULI(3'd7, 32'h00000001, 32'h7fffffff)
`STIMULI(3'd7, 32'h00000000, 32'h7fffffff)
`STIMULI(3'd7, 32'hffffffff, 32'h00000002)
`STIMULI(3'd7, 32'hfffffffe, 32'h00000002)
`STIMULI(3'd7, 32'h80000001, 32'h00000002)
`STIMULI(3'd7, 32'h80000000, 32'h00000002)
`STIMULI(3'd7, 32'h7fffffff, 32'h00000002)
`STIMULI(3'd7, 32'h00000002, 32'h00000002)
`STIMULI(3'd7, 32'h00000001, 32'h00000002)
`STIMULI(3'd7, 32'h00000000, 32'h00000002)
`STIMULI(3'd7, 32'hffffffff, 32'h00000001)
`STIMULI(3'd7, 32'hfffffffe, 32'h00000001)
`STIMULI(3'd7, 32'h80000001, 32'h00000001)
`STIMULI(3'd7, 32'h80000000, 32'h00000001)
`STIMULI(3'd7, 32'h7fffffff, 32'h00000001)
`STIMULI(3'd7, 32'h00000002, 32'h00000001)
`STIMULI(3'd7, 32'h00000001, 32'h00000001)
`STIMULI(3'd7, 32'h00000000, 32'h00000001)
`STIMULI(3'd7, 32'hffffffff, 32'h00000000)
`STIMULI(3'd7, 32'hfffffffe, 32'h00000000)
`STIMULI(3'd7, 32'h80000001, 32'h00000000)
`STIMULI(3'd7, 32'h80000000, 32'h00000000)
`STIMULI(3'd7, 32'h7fffffff, 32'h00000000)
`STIMULI(3'd7, 32'h00000002, 32'h00000000)
`STIMULI(3'd7, 32'h00000001, 32'h00000000)
`STIMULI(3'd7, 32'h00000000, 32'h00000000)
`STIMULI(3'd7, 32'h5ece7607, 32'h322e104d)
`STIMULI(3'd7, 32'hafbf9f22, 32'hb46c1093)
`STIMULI(3'd7, 32'hb63ab2dd, 32'hbc01362a)
`STIMULI(3'd7, 32'h2d57f6db, 32'h950928e4)
`STIMULI(3'd7, 32'h6e2f4677, 32'h5d1795fd)
`STIMULI(3'd7, 32'h49753977, 32'h2469f954)
`STIMULI(3'd7, 32'h1918cc27, 32'h76cd3052)
`STIMULI(3'd7, 32'h39732238, 32'h8748129f)
`STIMULI(3'd7, 32'h53e4c650, 32'h02e85baf)
`STIMULI(3'd7, 32'h2bb20bf3, 32'h6cfd9277)
`STIMULI(3'd7, 32'h79b58c02, 32'h65252e2c)
`STIMULI(3'd7, 32'h7445a516, 32'h4d9a5252)
`STIMULI(3'd7, 32'h680d89db, 32'h9ff7b10a)
`STIMULI(3'd7, 32'h3a97e4c9, 32'h61c315dd)
`STIMULI(3'd7, 32'h851cdf36, 32'haedd89e0)
`STIMULI(3'd7, 32'h2f5d682f, 32'h6d2a6911)
`STIMULI(3'd7, 32'h4ed53aea, 32'h69f54cf9)
`STIMULI(3'd7, 32'h4eed7eef, 32'h53f21a20)
`STIMULI(3'd7, 32'h98d2d6d9, 32'h7e4ae71e)
`STIMULI(3'd7, 32'h411c8331, 32'h67a811c3)
`STIMULI(3'd7, 32'h68403417, 32'h100a0220)
`STIMULI(3'd7, 32'hbb9a2be3, 32'h01130af0)
`STIMULI(3'd7, 32'h8e54e93f, 32'h7cb6af14)
`STIMULI(3'd7, 32'h68bb1cb3, 32'h76951d56)
`STIMULI(3'd7, 32'h8cc0b135, 32'h24554896)
`STIMULI(3'd7, 32'h77a82847, 32'h9b159a74)
`STIMULI(3'd7, 32'ha10bf7ab, 32'h606344fa)
`STIMULI(3'd7, 32'h11aab7ca, 32'hadcca8e0)
`STIMULI(3'd7, 32'h84b88d91, 32'h0952e011)
`STIMULI(3'd7, 32'h48e24354, 32'ha5c4853c)
`STIMULI(3'd7, 32'h69b6250c, 32'h5a8cfb1e)
`STIMULI(3'd7, 32'h53912e1c, 32'h6e6eb29d)
`STIMULI(3'd7, 32'h63dfdb30, 32'h9c737170)
`STIMULI(3'd7, 32'h943337d9, 32'h4d96003c)
`STIMULI(3'd7, 32'h77006c8e, 32'h67c465f5)
`STIMULI(3'd7, 32'hbc04b2d9, 32'h5ae047be)
`STIMULI(3'd7, 32'h8437d765, 32'h5037eab2)
`STIMULI(3'd7, 32'h287647fa, 32'h7b3843f3)
`STIMULI(3'd7, 32'hb7fc50a7, 32'h647afad3)
`STIMULI(3'd7, 32'h56188bb2, 32'hbc34280c)
`STIMULI(3'd7, 32'h34b2e585, 32'h7e8ed3ac)
`STIMULI(3'd7, 32'h376c6bff, 32'h6caf362c)
`STIMULI(3'd7, 32'h6309ce80, 32'h0d84f7b1)
`STIMULI(3'd7, 32'h28e35e38, 32'h17bcb405)
`STIMULI(3'd7, 32'h8c13cb5e, 32'h604fca38)
`STIMULI(3'd7, 32'h846bea32, 32'h6f1d99de)
`STIMULI(3'd7, 32'h6dd4c1e9, 32'h2d4f486a)
`STIMULI(3'd7, 32'h06da4de3, 32'h79e88d47)
`STIMULI(3'd7, 32'h0d9f12a2, 32'h0b463815)
`STIMULI(3'd7, 32'h69062725, 32'h7b73d48c)
`STIMULI(3'd7, 32'hb8958080, 32'h6fe07509)
`STIMULI(3'd7, 32'h755c61d3, 32'h46349322)
`STIMULI(3'd7, 32'h7b26ad1e, 32'h5e6288f9)
`STIMULI(3'd7, 32'h41a867ae, 32'h33bc2d9e)
`STIMULI(3'd7, 32'h4e42fe02, 32'hb704c982)
`STIMULI(3'd7, 32'h79f0c0c1, 32'h4969ab20)
`STIMULI(3'd7, 32'h9567527b, 32'h3b99286f)
`STIMULI(3'd7, 32'h7d25d8bf, 32'h63aa507d)
`STIMULI(3'd7, 32'h729df1f1, 32'h77169980)
`STIMULI(3'd7, 32'h2d13fb9d, 32'h0805446c)
`STIMULI(3'd7, 32'h32afc1ef, 32'h2a39d45c)
`STIMULI(3'd7, 32'h6baf94e9, 32'ha54db3e1)
`STIMULI(3'd7, 32'h21506ddc, 32'h98c39087)
`STIMULI(3'd7, 32'h2d52f84d, 32'h54002fcc)
`STIMULI(3'd7, 32'h42fd64e3, 32'h99028d37)
`STIMULI(3'd7, 32'h794de3ad, 32'h644dd2c0)
`STIMULI(3'd7, 32'hb1c61dbe, 32'h26a0dbfa)
`STIMULI(3'd7, 32'hb84e028c, 32'h74c382a1)
`STIMULI(3'd7, 32'h3fa36931, 32'hb19be639)
