/* =========================================
* Top module wrapper of an accelerator role
*
* Author: Yisong Chang (changyisong@ict.ac.cn)
* Date: 29/01/2021
* Version: v0.0.1
*===========================================
*/

`timescale 10 ns / 1 ns

module custom_role (
  /* accelerator source clock */
  input        role_clk,
  input        role_resetn,

  /* memory interface clock */
  input        role_to_mem_clk,
  input        role_to_mem_resetn,

  /* AXI4 master: 
  *  to SHELL DDR4 memory controller */
  output [39:0] axi_role_to_mem_araddr,
  output [1:0]  axi_role_to_mem_arburst,
  output [3:0]  axi_role_to_mem_arcache,
  output [7:0]  axi_role_to_mem_arlen,
  output [0:0]  axi_role_to_mem_arlock,
  output [2:0]  axi_role_to_mem_arprot,
  output [3:0]  axi_role_to_mem_arqos,
  input         axi_role_to_mem_arready,
  output [3:0]	axi_role_to_mem_arregion,
  output [2:0]	axi_role_to_mem_arsize,
  output        axi_role_to_mem_arvalid,
  output [39:0]	axi_role_to_mem_awaddr,
  output [1:0]	axi_role_to_mem_awburst,
  output [3:0]	axi_role_to_mem_awcache,
  output [7:0]	axi_role_to_mem_awlen,
  output [0:0]	axi_role_to_mem_awlock,
  output [2:0]	axi_role_to_mem_awprot,
  output [3:0]	axi_role_to_mem_awqos,
  input         axi_role_to_mem_awready,
  output [3:0]	axi_role_to_mem_awregion,
  output [2:0]	axi_role_to_mem_awsize,
  output        axi_role_to_mem_awvalid,
  output        axi_role_to_mem_bready,
  input [1:0]   axi_role_to_mem_bresp,
  input         axi_role_to_mem_bvalid,
  input [63:0] axi_role_to_mem_rdata,
  input         axi_role_to_mem_rlast,
  output        axi_role_to_mem_rready,
  input [1:0]   axi_role_to_mem_rresp,
  input         axi_role_to_mem_rvalid,
  output [63:0] axi_role_to_mem_wdata,
  output        axi_role_to_mem_wlast,
  input         axi_role_to_mem_wready,
  output [7:0]  axi_role_to_mem_wstrb,
  output        axi_role_to_mem_wvalid,

  /* AXI4-lite master: 
  *  to SHELL UART controller and etc. */
  output [31:0] axi_role_to_shell_araddr,
  output [2:0]  axi_role_to_shell_arprot,
  input         axi_role_to_shell_arready,
  output        axi_role_to_shell_arvalid,
  output [31:0] axi_role_to_shell_awaddr,
  output [2:0]  axi_role_to_shell_awprot,
  input         axi_role_to_shell_awready,
  output        axi_role_to_shell_awvalid,
  output        axi_role_to_shell_bready,
  input [1:0]   axi_role_to_shell_bresp,
  input         axi_role_to_shell_bvalid,
  input [31:0]  axi_role_to_shell_rdata,
  output        axi_role_to_shell_rready,
  input [1:0]   axi_role_to_shell_rresp,
  input         axi_role_to_shell_rvalid,
  output [31:0] axi_role_to_shell_wdata,
  input         axi_role_to_shell_wready,
  output [3:0]  axi_role_to_shell_wstrb,
  output        axi_role_to_shell_wvalid,

  /* AXI4-lite slave: 
  *  from SHELL to MMIO registers in role */
  input [19:0]  axi_shell_to_role_araddr,
  input [2:0]   axi_shell_to_role_arprot,
  output        axi_shell_to_role_arready,
  input         axi_shell_to_role_arvalid,
  input [19:0]  axi_shell_to_role_awaddr,
  input [2:0]   axi_shell_to_role_awprot,
  output        axi_shell_to_role_awready,
  input         axi_shell_to_role_awvalid,
  input         axi_shell_to_role_bready,
  output [1:0]  axi_shell_to_role_bresp,
  output        axi_shell_to_role_bvalid,
  output [31:0] axi_shell_to_role_rdata,
  input         axi_shell_to_role_rready,
  output [1:0]  axi_shell_to_role_rresp,
  output        axi_shell_to_role_rvalid,
  input [31:0]  axi_shell_to_role_wdata,
  output        axi_shell_to_role_wready,
  input [3:0]   axi_shell_to_role_wstrb,
  input         axi_shell_to_role_wvalid
);

 role_wrapper role_wrapper_i (
    .axi_role_to_mem_araddr     (axi_role_to_mem_araddr   ),
    .axi_role_to_mem_arburst    (axi_role_to_mem_arburst  ),
    .axi_role_to_mem_arcache    (axi_role_to_mem_arcache  ),
    .axi_role_to_mem_arlen      (axi_role_to_mem_arlen    ),
    .axi_role_to_mem_arlock     (axi_role_to_mem_arlock   ),
    .axi_role_to_mem_arprot     (axi_role_to_mem_arprot   ),
    .axi_role_to_mem_arqos      (axi_role_to_mem_arqos    ),
    .axi_role_to_mem_arready    (axi_role_to_mem_arready  ),
    .axi_role_to_mem_arregion   (axi_role_to_mem_arregion ),
    .axi_role_to_mem_arsize     (axi_role_to_mem_arsize   ),
    .axi_role_to_mem_arvalid    (axi_role_to_mem_arvalid  ),
    .axi_role_to_mem_awaddr     (axi_role_to_mem_awaddr   ),
    .axi_role_to_mem_awburst    (axi_role_to_mem_awburst  ),
    .axi_role_to_mem_awcache    (axi_role_to_mem_awcache  ),
    .axi_role_to_mem_awlen      (axi_role_to_mem_awlen    ),
    .axi_role_to_mem_awlock     (axi_role_to_mem_awlock   ),
    .axi_role_to_mem_awprot     (axi_role_to_mem_awprot   ),
    .axi_role_to_mem_awqos      (axi_role_to_mem_awqos    ),
    .axi_role_to_mem_awready    (axi_role_to_mem_awready  ),
    .axi_role_to_mem_awregion   (axi_role_to_mem_awregion ),
    .axi_role_to_mem_awsize     (axi_role_to_mem_awsize   ),
    .axi_role_to_mem_awvalid    (axi_role_to_mem_awvalid  ),
    .axi_role_to_mem_bready     (axi_role_to_mem_bready   ),
    .axi_role_to_mem_bresp      (axi_role_to_mem_bresp    ),
    .axi_role_to_mem_bvalid     (axi_role_to_mem_bvalid   ),
    .axi_role_to_mem_rdata      (axi_role_to_mem_rdata    ),
    .axi_role_to_mem_rlast      (axi_role_to_mem_rlast    ),
    .axi_role_to_mem_rready     (axi_role_to_mem_rready   ),
    .axi_role_to_mem_rresp      (axi_role_to_mem_rresp    ),
    .axi_role_to_mem_rvalid     (axi_role_to_mem_rvalid   ),
    .axi_role_to_mem_wdata      (axi_role_to_mem_wdata    ),
    .axi_role_to_mem_wlast      (axi_role_to_mem_wlast    ),
    .axi_role_to_mem_wready     (axi_role_to_mem_wready   ),
    .axi_role_to_mem_wstrb      (axi_role_to_mem_wstrb    ),
    .axi_role_to_mem_wvalid     (axi_role_to_mem_wvalid   ),
    .axi_role_to_shell_araddr   (axi_role_to_shell_araddr ),
    .axi_role_to_shell_arprot   (axi_role_to_shell_arprot ),
    .axi_role_to_shell_arready  (axi_role_to_shell_arready),
    .axi_role_to_shell_arvalid  (axi_role_to_shell_arvalid),
    .axi_role_to_shell_awaddr   (axi_role_to_shell_awaddr ),
    .axi_role_to_shell_awprot   (axi_role_to_shell_awprot ),
    .axi_role_to_shell_awready  (axi_role_to_shell_awready),
    .axi_role_to_shell_awvalid  (axi_role_to_shell_awvalid),
    .axi_role_to_shell_bready   (axi_role_to_shell_bready ),
    .axi_role_to_shell_bresp    (axi_role_to_shell_bresp  ),
    .axi_role_to_shell_bvalid   (axi_role_to_shell_bvalid ),
    .axi_role_to_shell_rdata    (axi_role_to_shell_rdata  ),
    .axi_role_to_shell_rready   (axi_role_to_shell_rready ),
    .axi_role_to_shell_rresp    (axi_role_to_shell_rresp  ),
    .axi_role_to_shell_rvalid   (axi_role_to_shell_rvalid ),
    .axi_role_to_shell_wdata    (axi_role_to_shell_wdata  ),
    .axi_role_to_shell_wready   (axi_role_to_shell_wready ),
    .axi_role_to_shell_wstrb    (axi_role_to_shell_wstrb  ),
    .axi_role_to_shell_wvalid   (axi_role_to_shell_wvalid ),
    .axi_shell_to_role_araddr   (axi_shell_to_role_araddr ),
    .axi_shell_to_role_arprot   (axi_shell_to_role_arprot ),
    .axi_shell_to_role_arready  (axi_shell_to_role_arready),
    .axi_shell_to_role_arvalid  (axi_shell_to_role_arvalid),
    .axi_shell_to_role_awaddr   (axi_shell_to_role_awaddr ),
    .axi_shell_to_role_awprot   (axi_shell_to_role_awprot ),
    .axi_shell_to_role_awready  (axi_shell_to_role_awready),
    .axi_shell_to_role_awvalid  (axi_shell_to_role_awvalid),
    .axi_shell_to_role_bready   (axi_shell_to_role_bready ),
    .axi_shell_to_role_bresp    (axi_shell_to_role_bresp  ),
    .axi_shell_to_role_bvalid   (axi_shell_to_role_bvalid ),
    .axi_shell_to_role_rdata    (axi_shell_to_role_rdata  ),
    .axi_shell_to_role_rready   (axi_shell_to_role_rready ),
    .axi_shell_to_role_rresp    (axi_shell_to_role_rresp  ),
    .axi_shell_to_role_rvalid   (axi_shell_to_role_rvalid ),
    .axi_shell_to_role_wdata    (axi_shell_to_role_wdata  ),
    .axi_shell_to_role_wready   (axi_shell_to_role_wready ),
    .axi_shell_to_role_wstrb    (axi_shell_to_role_wstrb  ),
    .axi_shell_to_role_wvalid   (axi_shell_to_role_wvalid ),
    .role_clk                   (role_clk),
    .role_resetn                (role_resetn),
    .role_to_mem_clk            (role_to_mem_clk),
    .role_to_mem_resetn         (role_to_mem_resetn)
 );
 
 endmodule
