`STIMULI(5'h01, 5'h00, 5'h01, 32'h12153524, 1'h1)
`STIMULI(5'h02, 5'h01, 5'h02, 32'h1158a1b8, 1'h1)
`STIMULI(5'h03, 5'h02, 5'h03, 32'h78fdc89a, 1'h1)
`STIMULI(5'h10, 5'h03, 5'h10, 32'hec789fbb, 1'h1)
`STIMULI(5'h08, 5'h10, 5'h08, 32'hcd8acd8a, 1'h1)
`STIMULI(5'h00, 5'h08, 5'h00, 32'hdec87ac4, 1'h1)
`STIMULI(5'h01, 5'h08, 5'h01, 32'h12153524, 1'h1)
`STIMULI(5'h02, 5'h01, 5'h02, 32'h1158a1b8, 1'h0)
`STIMULI(5'h03, 5'h02, 5'h03, 32'h78fdc89a, 1'h0)
`STIMULI(5'h10, 5'h03, 5'h10, 32'hec789fbb, 1'h0)
`STIMULI(5'h08, 5'h10, 5'h08, 32'hcd8acd8a, 1'h0)
`STIMULI(5'h00, 5'h08, 5'h00, 32'hdec87ac4, 1'h0)
`STIMULI(5'h08, 5'h01, 5'h01, 32'h12153524, 1'h1)
`STIMULI(5'h01, 5'h02, 5'h02, 32'h1158a1b8, 1'h1)
`STIMULI(5'h02, 5'h03, 5'h03, 32'h78fdc89a, 1'h1)
`STIMULI(5'h03, 5'h10, 5'h10, 32'hec789fbb, 1'h1)
`STIMULI(5'h10, 5'h08, 5'h08, 32'hcd8acd8a, 1'h1)
`STIMULI(5'h08, 5'h00, 5'h00, 32'hdec87ac4, 1'h1)
`STIMULI(5'h08, 5'h01, 5'h01, 32'h12153524, 1'h1)
`STIMULI(5'h01, 5'h02, 5'h02, 32'h1158a1b8, 1'h0)
`STIMULI(5'h02, 5'h03, 5'h03, 32'h78fdc89a, 1'h0)
`STIMULI(5'h03, 5'h10, 5'h10, 32'hec789fbb, 1'h0)
`STIMULI(5'h10, 5'h08, 5'h08, 32'hcd8acd8a, 1'h0)
`STIMULI(5'h08, 5'h00, 5'h00, 32'hdec87ac4, 1'h0)
`STIMULI(5'h0d, 5'h0d, 5'h03, 32'hb1f05663, 1'h1)
`STIMULI(5'h03, 5'h03, 5'h03, 32'hc780c01a, 1'h1)
`STIMULI(5'h08, 5'h08, 5'h0d, 32'hb78cacd7, 1'h1)
`STIMULI(5'h0d, 5'h0d, 5'h0d, 32'hcd8a14ca, 1'h1)
`STIMULI(5'h00, 5'h00, 5'h05, 32'h78da5442, 1'h1)
`STIMULI(5'h0d, 5'h0d, 5'h03, 32'hb1f05663, 1'h0)
`STIMULI(5'h03, 5'h03, 5'h03, 32'hc780c01a, 1'h0)
`STIMULI(5'h08, 5'h08, 5'h0d, 32'hb78cacd7, 1'h0)
`STIMULI(5'h0d, 5'h0d, 5'h0d, 32'hcd8a14ca, 1'h0)
`STIMULI(5'h00, 5'h00, 5'h05, 32'h78da5442, 1'h0)
`STIMULI(5'h01, 5'h01, 5'h01, 32'h0aec3515, 1'h1)
`STIMULI(5'h05, 5'h05, 5'h05, 32'ha18bee43, 1'h1)
`STIMULI(5'h08, 5'h08, 5'h08, 32'h1297cb25, 1'h1)
`STIMULI(5'h10, 5'h10, 5'h10, 32'had67e25a, 1'h1)
`STIMULI(5'h17, 5'h17, 5'h17, 32'h060a5d0c, 1'h1)
`STIMULI(5'h1f, 5'h1f, 5'h1f, 32'h60decbc1, 1'h1)
`STIMULI(5'h00, 5'h00, 5'h00, 32'h5b60e5b6, 1'h1)
`STIMULI(5'h01, 5'h01, 5'h01, 32'h0aec3515, 1'h0)
`STIMULI(5'h05, 5'h05, 5'h05, 32'ha18bee43, 1'h0)
`STIMULI(5'h08, 5'h08, 5'h08, 32'h1297cb25, 1'h0)
`STIMULI(5'h10, 5'h10, 5'h10, 32'had67e25a, 1'h0)
`STIMULI(5'h17, 5'h17, 5'h17, 32'h060a5d0c, 1'h0)
`STIMULI(5'h1f, 5'h1f, 5'h1f, 32'h60decbc1, 1'h0)
`STIMULI(5'h00, 5'h00, 5'h00, 32'h5b60e5b6, 1'h0)
`STIMULI(5'h15, 5'h00, 5'h17, 32'hae78585c, 1'h1)
`STIMULI(5'h12, 5'h03, 5'h03, 32'hb2c28465, 1'h1)
`STIMULI(5'h16, 5'h16, 5'h16, 32'h06d7cd0d, 1'h1)
`STIMULI(5'h0c, 5'h19, 5'h05, 32'h76d457ed, 1'h1)
`STIMULI(5'h05, 5'h0a, 5'h06, 32'he33724c6, 1'h1)
`STIMULI(5'h17, 5'h12, 5'h07, 32'h72aff7e5, 1'h1)
`STIMULI(5'h12, 5'h0e, 5'h08, 32'h47ecdb8f, 1'h1)
`STIMULI(5'h05, 5'h1c, 5'h09, 32'hf4007ae8, 1'h1)
`STIMULI(5'h0d, 5'h05, 5'h0a, 32'hde8e28bd, 1'h1)
`STIMULI(5'h0a, 5'h00, 5'h0b, 32'hb1ef6263, 1'h1)
`STIMULI(5'h0a, 5'h1d, 5'h0c, 32'h10642120, 1'h1)
`STIMULI(5'h13, 5'h0d, 5'h0d, 32'hcb203e96, 1'h1)
`STIMULI(5'h0b, 5'h15, 5'h0e, 32'ha9a7d653, 1'h1)
`STIMULI(5'h0e, 5'h1d, 5'h0f, 32'h81174a02, 1'h1)
`STIMULI(5'h03, 5'h0a, 5'h10, 32'he7c572cf, 1'h1)
`STIMULI(5'h1c, 5'h12, 5'h11, 32'he5730aca, 1'h1)
`STIMULI(5'h01, 5'h18, 5'h12, 32'h452e618a, 1'h1)
`STIMULI(5'h09, 5'h0b, 5'h13, 32'h3c20f378, 1'h1)
`STIMULI(5'h06, 5'h0e, 5'h14, 32'h5b0265b6, 1'h1)
`STIMULI(5'h0a, 5'h0b, 5'h15, 32'hde7502bc, 1'h1)
`STIMULI(5'h05, 5'h0f, 5'h16, 32'hb897be71, 1'h1)
`STIMULI(5'h1a, 5'h1e, 5'h17, 32'h9dcc603b, 1'h1)
`STIMULI(5'h11, 5'h19, 5'h18, 32'h0aaa4b15, 1'h1)
`STIMULI(5'h0c, 5'h1f, 5'h19, 32'h31230762, 1'h1)
`STIMULI(5'h18, 5'h17, 5'h1a, 32'h47b9a18f, 1'h1)
`STIMULI(5'h1c, 5'h1b, 5'h1b, 32'hcfc4569f, 1'h1)
`STIMULI(5'h09, 5'h10, 5'h1c, 32'h44de3789, 1'h1)
`STIMULI(5'h11, 5'h16, 5'h1d, 32'hebfec0d7, 1'h1)
`STIMULI(5'h02, 5'h08, 5'h1e, 32'h061d7f0c, 1'h1)
`STIMULI(5'h1d, 5'h12, 5'h1f, 32'hbb825a77, 1'h1)
`STIMULI(5'h0d, 5'h19, 5'h00, 32'hbf05007e, 1'h1)
`STIMULI(5'h13, 5'h05, 5'h01, 32'h0fd28f1f, 1'h1)
`STIMULI(5'h1b, 5'h09, 5'h02, 32'hbc148878, 1'h1)
`STIMULI(5'h0a, 5'h18, 5'h03, 32'h9ff2ae3f, 1'h1)
`STIMULI(5'h0e, 5'h1c, 5'h04, 32'hc33f3886, 1'h1)
`STIMULI(5'h06, 5'h13, 5'h05, 32'h7d3599fa, 1'h1)
`STIMULI(5'h0f, 5'h13, 5'h06, 32'hd18bb4a3, 1'h1)
`STIMULI(5'h04, 5'h17, 5'h07, 32'hafd8565f, 1'h1)
`STIMULI(5'h06, 5'h1a, 5'h08, 32'he59b36cb, 1'h1)
`STIMULI(5'h0d, 5'h1a, 5'h09, 32'h14cfc129, 1'h1)
`STIMULI(5'h15, 5'h1f, 5'h0a, 32'hb29fb665, 1'h1)
`STIMULI(5'h04, 5'h10, 5'h0b, 32'h3cf11979, 1'h1)
`STIMULI(5'h0b, 5'h0e, 5'h0c, 32'h15090b2a, 1'h1)
`STIMULI(5'h1a, 5'h1d, 5'h0d, 32'h6e5daddc, 1'h1)
`STIMULI(5'h16, 5'h0e, 5'h0e, 32'he1f102c3, 1'h1)
`STIMULI(5'h0a, 5'h16, 5'h0f, 32'hb3d97667, 1'h1)
`STIMULI(5'h19, 5'h18, 5'h10, 32'h9c0e8a38, 1'h1)
`STIMULI(5'h13, 5'h04, 5'h11, 32'h4a74bf94, 1'h1)
`STIMULI(5'h1b, 5'h0d, 5'h12, 32'hacb7ca59, 1'h1)
`STIMULI(5'h0d, 5'h16, 5'h13, 32'h6cb0b7d9, 1'h1)
`STIMULI(5'h16, 5'h15, 5'h14, 32'h653b49ca, 1'h0)
`STIMULI(5'h04, 5'h17, 5'h15, 32'ha3071a46, 1'h1)
`STIMULI(5'h14, 5'h08, 5'h16, 32'h34980769, 1'h1)
`STIMULI(5'h0d, 5'h07, 5'h17, 32'h147cd928, 1'h1)
`STIMULI(5'h08, 5'h1c, 5'h18, 32'h975c9c2e, 1'h1)
`STIMULI(5'h09, 5'h1c, 5'h19, 32'hfea7a6fd, 1'h1)
`STIMULI(5'h1a, 5'h1d, 5'h1a, 32'h43356786, 1'h1)
`STIMULI(5'h10, 5'h13, 5'h1b, 32'h334ea766, 1'h0)
`STIMULI(5'h1e, 5'h1a, 5'h1c, 32'h5d7199ba, 1'h1)
`STIMULI(5'h1a, 5'h19, 5'h1d, 32'h6a8e05d5, 1'h1)
`STIMULI(5'h16, 5'h00, 5'h1e, 32'h1b876137, 1'h0)
`STIMULI(5'h16, 5'h1d, 5'h1f, 32'h13259f26, 1'h1)
`STIMULI(5'h06, 5'h18, 5'h00, 32'h6e5f0fdc, 1'h1)
`STIMULI(5'h1b, 5'h0f, 5'h01, 32'h3f5a9b7e, 1'h0)
`STIMULI(5'h1a, 5'h01, 5'h02, 32'h3ced2b79, 1'h1)
`STIMULI(5'h01, 5'h06, 5'h03, 32'h0b940917, 1'h0)
`STIMULI(5'h15, 5'h15, 5'h04, 32'ha8639650, 1'h1)
`STIMULI(5'h01, 5'h05, 5'h05, 32'h949a8a29, 1'h0)
`STIMULI(5'h0b, 5'h13, 5'h06, 32'hcc01b498, 1'h1)
`STIMULI(5'h0a, 5'h0e, 5'h07, 32'hf622e6ec, 1'h1)
`STIMULI(5'h09, 5'h01, 5'h08, 32'hd44b80a8, 1'h0)
`STIMULI(5'h06, 5'h1f, 5'h09, 32'h070bb90e, 1'h1)
`STIMULI(5'h0a, 5'h0d, 5'h0a, 32'h152fb52a, 1'h0)
`STIMULI(5'h18, 5'h19, 5'h0b, 32'h4f75ff9e, 1'h0)
`STIMULI(5'h0a, 5'h13, 5'h0c, 32'h6464e3c8, 1'h0)
`STIMULI(5'h07, 5'h16, 5'h0d, 32'h35a0c96b, 1'h1)
`STIMULI(5'h04, 5'h19, 5'h0e, 32'h5d059dba, 1'h0)
`STIMULI(5'h14, 5'h1f, 5'h0f, 32'h492fd392, 1'h1)
`STIMULI(5'h1a, 5'h12, 5'h10, 32'hc3339086, 1'h1)
`STIMULI(5'h1d, 5'h04, 5'h11, 32'h19452132, 1'h1)
`STIMULI(5'h0a, 5'h09, 5'h12, 32'hf249a4e4, 1'h1)
`STIMULI(5'h0e, 5'h1b, 5'h13, 32'hd095a8a1, 1'h0)
`STIMULI(5'h0f, 5'h09, 5'h14, 32'h85e51e0b, 1'h0)
`STIMULI(5'h15, 5'h0f, 5'h15, 32'h1b60e536, 1'h0)
`STIMULI(5'h08, 5'h0e, 5'h16, 32'h35cdbf6b, 1'h0)
`STIMULI(5'h12, 5'h08, 5'h17, 32'h4df3819b, 1'h1)
`STIMULI(5'h0b, 5'h02, 5'h18, 32'h9684e02d, 1'h0)
`STIMULI(5'h0d, 5'h0c, 5'h19, 32'h8f1cf61e, 1'h1)
`STIMULI(5'h11, 5'h06, 5'h1a, 32'h0c039d18, 1'h1)
`STIMULI(5'h1b, 5'h18, 5'h1b, 32'ha0c02441, 1'h1)
`STIMULI(5'h16, 5'h1b, 5'h1c, 32'h29efe953, 1'h1)
`STIMULI(5'h04, 5'h13, 5'h1d, 32'hf166fae2, 1'h1)
`STIMULI(5'h12, 5'h18, 5'h1e, 32'hec50b4d8, 1'h0)
`STIMULI(5'h05, 5'h01, 5'h1f, 32'h9c811239, 1'h0)
`STIMULI(5'h01, 5'h08, 5'h00, 32'h15890f2b, 1'h1)
`STIMULI(5'h01, 5'h1f, 5'h01, 32'h13b55527, 1'h1)
`STIMULI(5'h18, 5'h16, 5'h02, 32'h82223a04, 1'h1)
`STIMULI(5'h12, 5'h16, 5'h03, 32'h0a6e9314, 1'h0)
`STIMULI(5'h15, 5'h0d, 5'h04, 32'hd8ace2b1, 1'h0)
`STIMULI(5'h15, 5'h0d, 5'h05, 32'h158b2b2b, 1'h0)
`STIMULI(5'h04, 5'h07, 5'h06, 32'h93c12227, 1'h0)
`STIMULI(5'h19, 5'h09, 5'h07, 32'hf3d7a6e7, 1'h0)
`STIMULI(5'h09, 5'h11, 5'h08, 32'h6de5bbdb, 1'h1)
`STIMULI(5'h0a, 5'h1a, 5'h09, 32'hd0bc5ea1, 1'h0)
`STIMULI(5'h03, 5'h1c, 5'h0a, 32'ha2e62045, 1'h0)
`STIMULI(5'h1e, 5'h08, 5'h0b, 32'hb9461472, 1'h1)
`STIMULI(5'h06, 5'h10, 5'h0c, 32'hb7dfaa6f, 1'h1)
`STIMULI(5'h00, 5'h08, 5'h0d, 32'h1c719738, 1'h0)
`STIMULI(5'h05, 5'h00, 5'h0e, 32'h7b0da9f6, 1'h0)
`STIMULI(5'h19, 5'h10, 5'h0f, 32'h3a625f74, 1'h0)
`STIMULI(5'h0a, 5'h02, 5'h10, 32'h1e1c873c, 1'h0)
`STIMULI(5'h01, 5'h17, 5'h11, 32'h0aec3515, 1'h0)
`STIMULI(5'h09, 5'h06, 5'h12, 32'ha18bee43, 1'h1)
`STIMULI(5'h01, 5'h0d, 5'h13, 32'h1297cb25, 1'h1)
`STIMULI(5'h07, 5'h0c, 5'h14, 32'had67e25a, 1'h1)
`STIMULI(5'h11, 5'h1b, 5'h15, 32'h060a5d0c, 1'h1)
`STIMULI(5'h17, 5'h1e, 5'h16, 32'h5b60e5b6, 1'h1)
`STIMULI(5'h15, 5'h00, 5'h17, 32'hae78585c, 1'h0)
`STIMULI(5'h12, 5'h14, 5'h18, 32'hd00b12a0, 1'h0)
`STIMULI(5'h0d, 5'h0b, 5'h19, 32'h6e8af5dd, 1'h1)
`STIMULI(5'h1e, 5'h1d, 5'h1a, 32'hbccc4279, 1'h1)
`STIMULI(5'h0f, 5'h03, 5'h1b, 32'hbde0d27b, 1'h1)
`STIMULI(5'h1d, 5'h11, 5'h1c, 32'h71c129e3, 1'h0)
`STIMULI(5'h15, 5'h00, 5'h1d, 32'h22119f44, 1'h0)
`STIMULI(5'h12, 5'h18, 5'h1e, 32'hf6a178ed, 1'h1)
`STIMULI(5'h12, 5'h04, 5'h1f, 32'h46dcb78d, 1'h1)
`STIMULI(5'h0c, 5'h10, 5'h00, 32'h236afd46, 1'h0)
`STIMULI(5'h0a, 5'h04, 5'h01, 32'h0beac117, 1'h1)
`STIMULI(5'h1c, 5'h00, 5'h02, 32'hd55bbcaa, 1'h1)
`STIMULI(5'h0b, 5'h06, 5'h03, 32'h5d4a4dba, 1'h0)
`STIMULI(5'h12, 5'h02, 5'h04, 32'h92831e25, 1'h1)
`STIMULI(5'h14, 5'h1d, 5'h05, 32'ha48f7c49, 1'h1)
`STIMULI(5'h1c, 5'h07, 5'h06, 32'h25f2034b, 1'h1)
`STIMULI(5'h19, 5'h14, 5'h07, 32'h433e9786, 1'h0)
`STIMULI(5'h0c, 5'h0c, 5'h08, 32'h6851e5d0, 1'h1)
`STIMULI(5'h0a, 5'h11, 5'h09, 32'h03e9b707, 1'h1)
`STIMULI(5'h0b, 5'h13, 5'h0a, 32'h746affe8, 1'h0)
`STIMULI(5'h03, 5'h04, 5'h0b, 32'h76295bec, 1'h0)
`STIMULI(5'h19, 5'h1f, 5'h0c, 32'h64e165c9, 1'h0)
`STIMULI(5'h07, 5'h1d, 5'h0d, 32'hea5814d4, 1'h0)
`STIMULI(5'h02, 5'h09, 5'h0e, 32'h583125b0, 1'h1)
`STIMULI(5'h00, 5'h1c, 5'h0f, 32'hecb91ad9, 1'h1)
`STIMULI(5'h03, 5'h0a, 5'h10, 32'h49b16f93, 1'h0)
`STIMULI(5'h1d, 5'h1a, 5'h11, 32'he471f8c8, 1'h0)
`STIMULI(5'h0b, 5'h19, 5'h12, 32'h4226a984, 1'h1)
`STIMULI(5'h12, 5'h19, 5'h13, 32'h897f1c12, 1'h1)
`STIMULI(5'h0e, 5'h17, 5'h14, 32'he82b96d0, 1'h1)
`STIMULI(5'h06, 5'h1b, 5'h15, 32'h6d8b87db, 1'h1)
`STIMULI(5'h0f, 5'h09, 5'h16, 32'h80797c00, 1'h1)
`STIMULI(5'h19, 5'h05, 5'h17, 32'h8653620c, 1'h0)
`STIMULI(5'h10, 5'h11, 5'h18, 32'h67d735cf, 1'h1)
`STIMULI(5'h17, 5'h0a, 5'h19, 32'hb4f9a469, 1'h1)
`STIMULI(5'h1b, 5'h04, 5'h1a, 32'hec3758d8, 1'h1)
`STIMULI(5'h17, 5'h06, 5'h1b, 32'h5c78b1b8, 1'h0)
`STIMULI(5'h17, 5'h15, 5'h1c, 32'h984d5a30, 1'h0)
`STIMULI(5'h07, 5'h16, 5'h1d, 32'h6a15f5d4, 1'h0)
`STIMULI(5'h0b, 5'h01, 5'h1e, 32'h74a1ade9, 1'h0)
`STIMULI(5'h00, 5'h02, 5'h1f, 32'h6d808bdb, 1'h0)
`STIMULI(5'h10, 5'h0f, 5'h00, 32'he2ecdac5, 1'h0)
`STIMULI(5'h0f, 5'h09, 5'h01, 32'hb302da66, 1'h0)
`STIMULI(5'h06, 5'h0f, 5'h02, 32'h7c41aff8, 1'h1)
`STIMULI(5'h15, 5'h0e, 5'h03, 32'h70ef37e1, 1'h1)
`STIMULI(5'h05, 5'h08, 5'h04, 32'h304e4d60, 1'h1)
`STIMULI(5'h09, 5'h01, 5'h05, 32'h322f7d64, 1'h1)
`STIMULI(5'h0e, 5'h01, 5'h06, 32'hbbbc5277, 1'h1)
`STIMULI(5'h08, 5'h10, 5'h07, 32'h6a9fb9d5, 1'h0)
`STIMULI(5'h0f, 5'h11, 5'h08, 32'hd57800aa, 1'h1)
`STIMULI(5'h0e, 5'h02, 5'h09, 32'hbe9bbc7d, 1'h1)
`STIMULI(5'h09, 5'h0f, 5'h0a, 32'h1e664d3c, 1'h0)
`STIMULI(5'h0f, 5'h0a, 5'h0b, 32'hade7d05b, 1'h0)
`STIMULI(5'h13, 5'h13, 5'h0c, 32'h5cd20db9, 1'h1)
`STIMULI(5'h11, 5'h17, 5'h0d, 32'h32dc4165, 1'h1)
`STIMULI(5'h1a, 5'h11, 5'h0e, 32'hcc981099, 1'h0)
`STIMULI(5'h04, 5'h0a, 5'h0f, 32'h317c0762, 1'h1)
`STIMULI(5'h19, 5'h05, 5'h10, 32'hbeda447d, 1'h1)
`STIMULI(5'h09, 5'h01, 5'h11, 32'h76de6bed, 1'h1)
`STIMULI(5'h1b, 5'h0d, 5'h12, 32'h57c1d1af, 1'h1)
`STIMULI(5'h06, 5'h02, 5'h13, 32'h38139f70, 1'h0)
`STIMULI(5'h0a, 5'h1c, 5'h14, 32'h5e983dbd, 1'h0)
`STIMULI(5'h1b, 5'h05, 5'h15, 32'ha86c5e50, 1'h0)
`STIMULI(5'h16, 5'h1c, 5'h16, 32'hbc3f8478, 1'h1)
`STIMULI(5'h19, 5'h08, 5'h17, 32'h11cc9b23, 1'h0)
`STIMULI(5'h0e, 5'h13, 5'h18, 32'hddd146bb, 1'h0)
`STIMULI(5'h0e, 5'h14, 5'h19, 32'h0671030c, 1'h0)
`STIMULI(5'h19, 5'h13, 5'h1a, 32'hacecdc59, 1'h1)
`STIMULI(5'h15, 5'h0c, 5'h1b, 32'h7a4fbff4, 1'h1)
`STIMULI(5'h02, 5'h15, 5'h1c, 32'h9cfc7a39, 1'h0)
`STIMULI(5'h0e, 5'h02, 5'h1d, 32'h02fbf905, 1'h0)
`STIMULI(5'h08, 5'h0d, 5'h1e, 32'h5c7951b8, 1'h1)
`STIMULI(5'h08, 5'h10, 5'h1f, 32'hd7b48eaf, 1'h0)
`STIMULI(5'h0c, 5'h1b, 5'h00, 32'h7af6abf5, 1'h0)
`STIMULI(5'h05, 5'h0d, 5'h01, 32'ha005a640, 1'h0)
`STIMULI(5'h0d, 5'h09, 5'h02, 32'hb87c1070, 1'h1)
`STIMULI(5'h10, 5'h00, 5'h03, 32'h5e2551bc, 1'h0)
`STIMULI(5'h01, 5'h0d, 5'h04, 32'h28766950, 1'h0)
`STIMULI(5'h15, 5'h1d, 5'h05, 32'hfaf32ef5, 1'h1)
`STIMULI(5'h0a, 5'h1c, 5'h06, 32'hca481294, 1'h0)
`STIMULI(5'h1e, 5'h1a, 5'h07, 32'hdc4308b8, 1'h1)
`STIMULI(5'h07, 5'h13, 5'h08, 32'h23400b46, 1'h1)
`STIMULI(5'h17, 5'h05, 5'h09, 32'haada7455, 1'h1)
`STIMULI(5'h19, 5'h06, 5'h0a, 32'hb1800a63, 1'h1)
`STIMULI(5'h1e, 5'h10, 5'h0b, 32'hb4497668, 1'h1)
`STIMULI(5'h1c, 5'h19, 5'h0c, 32'h2d19a55a, 1'h0)
`STIMULI(5'h10, 5'h0f, 5'h0d, 32'h55861fab, 1'h0)
`STIMULI(5'h05, 5'h0d, 5'h0e, 32'h6c6a6dd8, 1'h0)
`STIMULI(5'h1c, 5'h1c, 5'h0f, 32'h45f3238b, 1'h1)
`STIMULI(5'h19, 5'h05, 5'h10, 32'hd27f0aa4, 1'h0)
`STIMULI(5'h13, 5'h18, 5'h11, 32'h9f398e3e, 1'h0)
`STIMULI(5'h1c, 5'h06, 5'h12, 32'h62056bc4, 1'h1)
`STIMULI(5'h18, 5'h05, 5'h13, 32'hcd1d509a, 1'h1)
`STIMULI(5'h1a, 5'h03, 5'h14, 32'h5515d1aa, 1'h0)
`STIMULI(5'h0c, 5'h09, 5'h15, 32'h5934e9b2, 1'h0)
`STIMULI(5'h0b, 5'h18, 5'h16, 32'h61dafdc3, 1'h0)
`STIMULI(5'h09, 5'h0f, 5'h17, 32'h792c03f2, 1'h1)
`STIMULI(5'h0d, 5'h08, 5'h18, 32'h0de14b1b, 1'h1)
`STIMULI(5'h0f, 5'h0b, 5'h19, 32'h92f91225, 1'h0)
`STIMULI(5'h00, 5'h1d, 5'h1a, 32'h8d94d21b, 1'h0)
`STIMULI(5'h04, 5'h17, 5'h1b, 32'h412dfd82, 1'h0)
`STIMULI(5'h12, 5'h19, 5'h1c, 32'h1b368b36, 1'h1)
`STIMULI(5'h16, 5'h0a, 5'h1d, 32'hf24baee4, 1'h1)
`STIMULI(5'h0e, 5'h0c, 5'h1e, 32'h605065c0, 1'h0)
`STIMULI(5'h1b, 5'h1c, 5'h1f, 32'hb8c0c271, 1'h0)
`STIMULI(5'h17, 5'h01, 5'h00, 32'hee7068dc, 1'h0)
`STIMULI(5'h15, 5'h09, 5'h01, 32'h75fb21eb, 1'h1)
`STIMULI(5'h1f, 5'h10, 5'h02, 32'hc7b2e28f, 1'h0)
`STIMULI(5'h16, 5'h02, 5'h03, 32'he9b49ad3, 1'h0)
`STIMULI(5'h11, 5'h17, 5'h04, 32'h0d63751a, 1'h1)
`STIMULI(5'h11, 5'h0d, 5'h05, 32'h87628e0e, 1'h0)
`STIMULI(5'h1c, 5'h18, 5'h06, 32'h02bd4305, 1'h0)
`STIMULI(5'h0a, 5'h05, 5'h07, 32'hf67088ec, 1'h0)
`STIMULI(5'h03, 5'h1e, 5'h08, 32'h1b920537, 1'h1)
`STIMULI(5'h1e, 5'h08, 5'h09, 32'hfeaddcfd, 1'h0)
`STIMULI(5'h10, 5'h06, 5'h0a, 32'hba603874, 1'h1)
`STIMULI(5'h08, 5'h05, 5'h0b, 32'h09164d12, 1'h1)
`STIMULI(5'h16, 5'h13, 5'h0c, 32'hff202efe, 1'h0)
`STIMULI(5'h0b, 5'h17, 5'h0d, 32'h7dddabfb, 1'h0)
`STIMULI(5'h14, 5'h0a, 5'h0e, 32'h87d0360f, 1'h0)
`STIMULI(5'h14, 5'h0b, 5'h0f, 32'hd3666ea6, 1'h0)
`STIMULI(5'h04, 5'h14, 5'h10, 32'hb587c26b, 1'h1)
`STIMULI(5'h01, 5'h05, 5'h11, 32'h468b618d, 1'h0)
`STIMULI(5'h09, 5'h00, 5'h12, 32'hdc9974b9, 1'h0)
`STIMULI(5'h1c, 5'h17, 5'h13, 32'ha3643246, 1'h0)
`STIMULI(5'h13, 5'h0e, 5'h14, 32'h2c0c5558, 1'h0)
`STIMULI(5'h10, 5'h10, 5'h15, 32'h6e6d23dc, 1'h1)
`STIMULI(5'h03, 5'h18, 5'h16, 32'h0073e500, 1'h1)
`STIMULI(5'h13, 5'h18, 5'h17, 32'hd0b99aa1, 1'h1)
`STIMULI(5'h07, 5'h1a, 5'h18, 32'h2fef3d5f, 1'h0)
`STIMULI(5'h10, 5'h0b, 5'h19, 32'h1699d12d, 1'h1)
`STIMULI(5'h12, 5'h0c, 5'h1a, 32'h98d73831, 1'h1)
`STIMULI(5'h15, 5'h00, 5'h1b, 32'h06db6b0d, 1'h1)
`STIMULI(5'h14, 5'h00, 5'h1c, 32'h4a638d94, 1'h0)
`STIMULI(5'h03, 5'h0d, 5'h1d, 32'h098d1513, 1'h0)
`STIMULI(5'h18, 5'h07, 5'h1e, 32'hee4ee6dc, 1'h1)
`STIMULI(5'h03, 5'h0b, 5'h1f, 32'hafed265f, 1'h1)
`STIMULI(5'h02, 5'h09, 5'h00, 32'h1c421738, 1'h1)
`STIMULI(5'h02, 5'h0e, 5'h01, 32'he3eb4cc7, 1'h1)
`STIMULI(5'h04, 5'h1b, 5'h02, 32'he38e22c7, 1'h1)
`STIMULI(5'h15, 5'h15, 5'h03, 32'h84651408, 1'h0)
`STIMULI(5'h18, 5'h02, 5'h04, 32'h8d7d721a, 1'h1)
`STIMULI(5'h10, 5'h03, 5'h05, 32'hac05a058, 1'h1)
`STIMULI(5'h05, 5'h0a, 5'h06, 32'h5243e3a4, 1'h0)
`STIMULI(5'h14, 5'h1b, 5'h07, 32'h03703906, 1'h0)
`STIMULI(5'h08, 5'h17, 5'h08, 32'he455f0c8, 1'h0)
`STIMULI(5'h15, 5'h11, 5'h09, 32'h7c1df3f8, 1'h0)
`STIMULI(5'h1b, 5'h15, 5'h0a, 32'h41aed583, 1'h1)
`STIMULI(5'h1b, 5'h0f, 5'h0b, 32'h581653b0, 1'h1)
`STIMULI(5'h18, 5'h1d, 5'h0c, 32'h984da630, 1'h0)
`STIMULI(5'h01, 5'h19, 5'h0d, 32'ha36ae846, 1'h0)
`STIMULI(5'h0f, 5'h0b, 5'h0e, 32'h2af17355, 1'h1)
`STIMULI(5'h13, 5'h08, 5'h0f, 32'hef1deade, 1'h0)
`STIMULI(5'h18, 5'h15, 5'h10, 32'h74dc69e9, 1'h0)
`STIMULI(5'h14, 5'h04, 5'h11, 32'h61dbe5c3, 1'h1)
`STIMULI(5'h16, 5'h0f, 5'h12, 32'h3f25ef7e, 1'h0)
`STIMULI(5'h00, 5'h02, 5'h13, 32'hc1b04483, 1'h0)
`STIMULI(5'h05, 5'h17, 5'h14, 32'h5fe3cbbf, 1'h1)
`STIMULI(5'h15, 5'h18, 5'h15, 32'h229d0b45, 1'h0)
`STIMULI(5'h0c, 5'h10, 5'h16, 32'h63323bc6, 1'h0)
`STIMULI(5'h1c, 5'h1c, 5'h17, 32'h18bd6331, 1'h1)
`STIMULI(5'h0e, 5'h09, 5'h18, 32'hd7e31eaf, 1'h1)
`STIMULI(5'h1e, 5'h05, 5'h19, 32'hd95b40b2, 1'h1)
`STIMULI(5'h08, 5'h02, 5'h1a, 32'h555c0faa, 1'h0)
`STIMULI(5'h13, 5'h1a, 5'h1b, 32'h4d20099a, 1'h0)
`STIMULI(5'h0b, 5'h02, 5'h1c, 32'hfdeb7cfb, 1'h0)
`STIMULI(5'h11, 5'h1e, 5'h1d, 32'he64828cc, 1'h1)
`STIMULI(5'h1b, 5'h1f, 5'h1e, 32'h309cdb61, 1'h0)
`STIMULI(5'h00, 5'h19, 5'h1f, 32'hc881bc91, 1'h0)
`STIMULI(5'h14, 5'h11, 5'h00, 32'hbf53b47e, 1'h1)
`STIMULI(5'h07, 5'h04, 5'h01, 32'ha4de2849, 1'h0)
`STIMULI(5'h1b, 5'h19, 5'h02, 32'h41b5d583, 1'h0)
`STIMULI(5'h17, 5'h11, 5'h03, 32'h4afebf95, 1'h0)
`STIMULI(5'h0f, 5'h04, 5'h04, 32'h732c5fe6, 1'h0)
`STIMULI(5'h1c, 5'h0b, 5'h05, 32'h89646012, 1'h1)
`STIMULI(5'h1f, 5'h02, 5'h06, 32'he203f0c4, 1'h0)
`STIMULI(5'h1a, 5'h00, 5'h07, 32'h398a1973, 1'h0)
`STIMULI(5'h14, 5'h1b, 5'h08, 32'hff73cafe, 1'h0)
`STIMULI(5'h02, 5'h1f, 5'h09, 32'h7132bbe2, 1'h1)
`STIMULI(5'h1f, 5'h10, 5'h0a, 32'hcc13e298, 1'h1)
`STIMULI(5'h1d, 5'h0b, 5'h0b, 32'h791189f2, 1'h0)
`STIMULI(5'h14, 5'h09, 5'h0c, 32'h5a0a0fb4, 1'h1)
`STIMULI(5'h0c, 5'h15, 5'h0d, 32'h89b5d413, 1'h1)
`STIMULI(5'h15, 5'h0f, 5'h0e, 32'h1df61f3b, 1'h1)
`STIMULI(5'h15, 5'h1c, 5'h0f, 32'h1a619934, 1'h1)
`STIMULI(5'h07, 5'h01, 5'h10, 32'hf964fef2, 1'h0)
`STIMULI(5'h01, 5'h09, 5'h11, 32'hf23316e4, 1'h1)
`STIMULI(5'h0d, 5'h1f, 5'h12, 32'hfd52d8fa, 1'h1)
`STIMULI(5'h08, 5'h0b, 5'h13, 32'hdac986b5, 1'h1)
`STIMULI(5'h17, 5'h0e, 5'h14, 32'h89042e12, 1'h0)
`STIMULI(5'h00, 5'h1a, 5'h15, 32'hfc4ca4f8, 1'h0)
`STIMULI(5'h0c, 5'h0a, 5'h16, 32'h913e0222, 1'h1)
`STIMULI(5'h1e, 5'h09, 5'h17, 32'h3d7f5b7a, 1'h0)
`STIMULI(5'h0b, 5'h0e, 5'h18, 32'hf5a4f2eb, 1'h0)
`STIMULI(5'h1c, 5'h05, 5'h19, 32'haf455e5e, 1'h1)
`STIMULI(5'h12, 5'h17, 5'h1a, 32'hc5cb548b, 1'h1)
`STIMULI(5'h01, 5'h0e, 5'h1b, 32'hc1c3d683, 1'h0)
`STIMULI(5'h15, 5'h0d, 5'h1c, 32'ha5365c4a, 1'h0)
`STIMULI(5'h14, 5'h0c, 5'h1d, 32'hf204eee4, 1'h1)
`STIMULI(5'h03, 5'h0c, 5'h1e, 32'h0d623f1a, 1'h0)
`STIMULI(5'h0d, 5'h1c, 5'h1f, 32'h79c681f3, 1'h0)
`STIMULI(5'h0c, 5'h0f, 5'h00, 32'h6e8d45dd, 1'h1)
`STIMULI(5'h18, 5'h0b, 5'h01, 32'h7fdbb3ff, 1'h0)
`STIMULI(5'h1b, 5'h13, 5'h02, 32'h13d1f727, 1'h1)
`STIMULI(5'h1b, 5'h06, 5'h03, 32'h06499b0c, 1'h1)
`STIMULI(5'h0a, 5'h0a, 5'h04, 32'ha4d83a49, 1'h0)
`STIMULI(5'h16, 5'h09, 5'h05, 32'h8c06d218, 1'h1)
`STIMULI(5'h1d, 5'h06, 5'h06, 32'h1725712e, 1'h0)
`STIMULI(5'h15, 5'h0f, 5'h07, 32'hbb062876, 1'h1)
`STIMULI(5'h1b, 5'h1c, 5'h08, 32'h4ad39595, 1'h0)
`STIMULI(5'h09, 5'h09, 5'h09, 32'hb7f4306f, 1'h0)
`STIMULI(5'h1a, 5'h0d, 5'h0a, 32'h5a3761b4, 1'h1)
`STIMULI(5'h0d, 5'h10, 5'h0b, 32'h6fcff1df, 1'h0)
`STIMULI(5'h11, 5'h04, 5'h0c, 32'h41bd6783, 1'h0)
`STIMULI(5'h19, 5'h06, 5'h0d, 32'hc0467280, 1'h0)
`STIMULI(5'h1f, 5'h09, 5'h0e, 32'he5063aca, 1'h1)
`STIMULI(5'h10, 5'h09, 5'h0f, 32'h42797584, 1'h1)
`STIMULI(5'h1e, 5'h0c, 5'h10, 32'h08098510, 1'h1)
`STIMULI(5'h17, 5'h01, 5'h11, 32'h0498fb09, 1'h1)
`STIMULI(5'h11, 5'h13, 5'h12, 32'h86c8320d, 1'h1)
`STIMULI(5'h0f, 5'h0e, 5'h13, 32'h4d77f99a, 1'h0)
`STIMULI(5'h06, 5'h1d, 5'h14, 32'h5bd583b7, 1'h1)
`STIMULI(5'h0f, 5'h04, 5'h15, 32'hce03ec9c, 1'h1)
`STIMULI(5'h02, 5'h09, 5'h16, 32'hcdbf3a9b, 1'h1)
`STIMULI(5'h0d, 5'h06, 5'h17, 32'h1747832e, 1'h0)
`STIMULI(5'h00, 5'h17, 5'h18, 32'hd51cb4aa, 1'h0)
`STIMULI(5'h08, 5'h0d, 5'h19, 32'hf8602ef0, 1'h0)
`STIMULI(5'h1b, 5'h1f, 5'h1a, 32'h68cd09d1, 1'h0)
`STIMULI(5'h18, 5'h1f, 5'h1b, 32'h3e8ed57d, 1'h0)
`STIMULI(5'h06, 5'h09, 5'h1c, 32'h4bac2f97, 1'h0)
`STIMULI(5'h17, 5'h1d, 5'h1d, 32'h624b63c4, 1'h1)
`STIMULI(5'h13, 5'h1f, 5'h1e, 32'h26c7134d, 1'h1)
`STIMULI(5'h19, 5'h00, 5'h1f, 32'ha703744e, 1'h1)
`STIMULI(5'h01, 5'h11, 5'h00, 32'h9cd6c239, 1'h1)
`STIMULI(5'h1e, 5'h1d, 5'h01, 32'h47ebef8f, 1'h1)
`STIMULI(5'h13, 5'h09, 5'h02, 32'h878a880f, 1'h1)
`STIMULI(5'h1a, 5'h1c, 5'h03, 32'h2b0da556, 1'h1)
`STIMULI(5'h13, 5'h1a, 5'h04, 32'h24e90749, 1'h0)
`STIMULI(5'h18, 5'h19, 5'h05, 32'h6c74f5d8, 1'h1)
`STIMULI(5'h09, 5'h16, 5'h06, 32'h92d06025, 1'h1)
`STIMULI(5'h13, 5'h1a, 5'h07, 32'h962c682c, 1'h1)
`STIMULI(5'h0c, 5'h08, 5'h08, 32'h005d5100, 1'h1)
`STIMULI(5'h00, 5'h1d, 5'h09, 32'hb66a586c, 1'h1)
`STIMULI(5'h00, 5'h1a, 5'h0a, 32'h68c14fd1, 1'h1)
`STIMULI(5'h00, 5'h0c, 5'h0b, 32'h6c1987d8, 1'h1)
`STIMULI(5'h11, 5'h11, 5'h0c, 32'he8cfb0d1, 1'h1)
`STIMULI(5'h13, 5'h1e, 5'h0d, 32'ha2a4be45, 1'h0)
`STIMULI(5'h1c, 5'h08, 5'h0e, 32'hc049c680, 1'h0)
`STIMULI(5'h11, 5'h07, 5'h0f, 32'hc0ad8081, 1'h1)
`STIMULI(5'h1f, 5'h00, 5'h10, 32'h41b1fd83, 1'h1)
`STIMULI(5'h1e, 5'h11, 5'h11, 32'hb2158c64, 1'h0)
`STIMULI(5'h1e, 5'h08, 5'h12, 32'h472dfb8e, 1'h0)
`STIMULI(5'h0a, 5'h1f, 5'h13, 32'h24839b49, 1'h0)
`STIMULI(5'h09, 5'h05, 5'h14, 32'ha8bfc851, 1'h0)
`STIMULI(5'h18, 5'h1e, 5'h15, 32'hb64ae66c, 1'h1)
`STIMULI(5'h03, 5'h07, 5'h16, 32'h97dde22f, 1'h0)
`STIMULI(5'h14, 5'h12, 5'h17, 32'h6a5ddbd4, 1'h0)
`STIMULI(5'h06, 5'h0f, 5'h18, 32'h1e32673c, 1'h0)
`STIMULI(5'h17, 5'h16, 5'h19, 32'ha0b3ae41, 1'h0)
`STIMULI(5'h02, 5'h03, 5'h1a, 32'h39092f72, 1'h0)
`STIMULI(5'h0b, 5'h08, 5'h1b, 32'hc9490292, 1'h0)
`STIMULI(5'h0b, 5'h15, 5'h1c, 32'h98b4ee31, 1'h1)
`STIMULI(5'h1e, 5'h0d, 5'h1d, 32'h38a38971, 1'h0)
`STIMULI(5'h08, 5'h02, 5'h1e, 32'hdaf356b5, 1'h0)
`STIMULI(5'h10, 5'h0c, 5'h1f, 32'h9f80983f, 1'h1)
`STIMULI(5'h05, 5'h1e, 5'h00, 32'h99183032, 1'h0)
`STIMULI(5'h1d, 5'h0a, 5'h01, 32'hdc16d8b8, 1'h0)
`STIMULI(5'h09, 5'h11, 5'h02, 32'hc6878a8d, 1'h0)
`STIMULI(5'h05, 5'h14, 5'h03, 32'hda12deb4, 1'h0)
`STIMULI(5'h0d, 5'h11, 5'h04, 32'h11c6c523, 1'h1)
`STIMULI(5'h14, 5'h0e, 5'h05, 32'h2f36c55e, 1'h1)
`STIMULI(5'h04, 5'h08, 5'h06, 32'h322cc164, 1'h1)
`STIMULI(5'h1b, 5'h0d, 5'h07, 32'hc544d88a, 1'h1)
`STIMULI(5'h0b, 5'h03, 5'h08, 32'hb5f8fa6b, 1'h1)
`STIMULI(5'h19, 5'h02, 5'h09, 32'h5e9d2fbd, 1'h0)
`STIMULI(5'h1f, 5'h1d, 5'h0a, 32'hf059ace0, 1'h1)
`STIMULI(5'h06, 5'h05, 5'h0b, 32'hc9b64c93, 1'h1)
`STIMULI(5'h0c, 5'h0b, 5'h0c, 32'h84a8e809, 1'h1)
`STIMULI(5'h17, 5'h05, 5'h0d, 32'h5858bdb0, 1'h0)
`STIMULI(5'h16, 5'h0f, 5'h0e, 32'habe8c057, 1'h1)
`STIMULI(5'h1d, 5'h07, 5'h0f, 32'h5a45bdb4, 1'h0)
`STIMULI(5'h06, 5'h1e, 5'h10, 32'h23466346, 1'h0)
`STIMULI(5'h14, 5'h14, 5'h11, 32'h1fb0d13f, 1'h1)
`STIMULI(5'h06, 5'h10, 5'h12, 32'ha62c344c, 1'h1)
`STIMULI(5'h06, 5'h0a, 5'h13, 32'h16b46d2d, 1'h0)
`STIMULI(5'h0f, 5'h00, 5'h14, 32'h5c2afdb8, 1'h1)
`STIMULI(5'h09, 5'h08, 5'h15, 32'h1fa98f3f, 1'h0)
`STIMULI(5'h1e, 5'h18, 5'h16, 32'haac1fa55, 1'h0)
`STIMULI(5'h16, 5'h05, 5'h17, 32'he70a62ce, 1'h1)
`STIMULI(5'h0f, 5'h15, 5'h18, 32'hd4ce0aa9, 1'h0)
`STIMULI(5'h16, 5'h15, 5'h19, 32'h2047dd40, 1'h0)
`STIMULI(5'h01, 5'h05, 5'h1a, 32'had27c45a, 1'h0)
`STIMULI(5'h04, 5'h19, 5'h1b, 32'h93ba6027, 1'h0)
`STIMULI(5'h08, 5'h09, 5'h1c, 32'hcfb89e9f, 1'h1)
`STIMULI(5'h05, 5'h13, 5'h1d, 32'h42955d85, 1'h1)
`STIMULI(5'h16, 5'h14, 5'h1e, 32'h440f0988, 1'h1)
`STIMULI(5'h11, 5'h1b, 5'h1f, 32'h1e85ed3d, 1'h1)
`STIMULI(5'h1d, 5'h14, 5'h00, 32'h8e39901c, 1'h0)
`STIMULI(5'h0f, 5'h19, 5'h01, 32'h2764754e, 1'h1)
`STIMULI(5'h1e, 5'h1d, 5'h02, 32'hf670fcec, 1'h1)
`STIMULI(5'h03, 5'h04, 5'h03, 32'he02148c0, 1'h1)
`STIMULI(5'h11, 5'h04, 5'h04, 32'ha5d9704b, 1'h1)
`STIMULI(5'h13, 5'h13, 5'h05, 32'h24d44749, 1'h1)
`STIMULI(5'h08, 5'h0a, 5'h06, 32'h0e62911c, 1'h1)
`STIMULI(5'h0e, 5'h0c, 5'h07, 32'h2e97795d, 1'h1)
`STIMULI(5'h18, 5'h0a, 5'h08, 32'h5d8e95bb, 1'h0)
`STIMULI(5'h1e, 5'h16, 5'h09, 32'h2e94b75d, 1'h1)
`STIMULI(5'h1b, 5'h14, 5'h0a, 32'h65a879cb, 1'h0)
`STIMULI(5'h04, 5'h19, 5'h0b, 32'h106e4320, 1'h1)
`STIMULI(5'h12, 5'h05, 5'h0c, 32'he6b110cd, 1'h0)
`STIMULI(5'h1e, 5'h1d, 5'h0d, 32'hd4ea6aa9, 1'h0)
`STIMULI(5'h0b, 5'h1b, 5'h0e, 32'h600b2dc0, 1'h1)
`STIMULI(5'h12, 5'h13, 5'h0f, 32'h408a2981, 1'h0)
`STIMULI(5'h08, 5'h01, 5'h10, 32'h05aeb90b, 1'h0)
`STIMULI(5'h0f, 5'h00, 5'h11, 32'h7e72c5fc, 1'h0)
`STIMULI(5'h15, 5'h19, 5'h12, 32'h076adf0e, 1'h0)
`STIMULI(5'h07, 5'h14, 5'h13, 32'h86d26e0d, 1'h0)
`STIMULI(5'h1f, 5'h1f, 5'h14, 32'h7e7f21fc, 1'h1)
`STIMULI(5'h08, 5'h1a, 5'h15, 32'hc0a7e881, 1'h0)
`STIMULI(5'h19, 5'h06, 5'h16, 32'hfd9380fb, 1'h0)
`STIMULI(5'h0f, 5'h0d, 5'h17, 32'h29951b53, 1'h0)
`STIMULI(5'h04, 5'h01, 5'h18, 32'h58d79db1, 1'h0)
`STIMULI(5'h08, 5'h14, 5'h19, 32'h7b24bdf6, 1'h0)
`STIMULI(5'h0a, 5'h1e, 5'h1a, 32'hb7d0ca6f, 1'h0)
`STIMULI(5'h06, 5'h1d, 5'h1b, 32'hfbaaeef7, 1'h1)
`STIMULI(5'h1a, 5'h14, 5'h1c, 32'hd01f40a0, 1'h0)
`STIMULI(5'h00, 5'h1c, 5'h1d, 32'h19a8e333, 1'h1)
`STIMULI(5'h09, 5'h0f, 5'h1e, 32'h38422d70, 1'h0)
`STIMULI(5'h17, 5'h03, 5'h1f, 32'h4b5b7196, 1'h0)
`STIMULI(5'h0a, 5'h0a, 5'h00, 32'h8322de06, 1'h1)
`STIMULI(5'h08, 5'h0d, 5'h01, 32'h20dcbf41, 1'h0)
`STIMULI(5'h08, 5'h13, 5'h02, 32'h38eedd71, 1'h1)
`STIMULI(5'h15, 5'h1e, 5'h03, 32'hb600e26c, 1'h1)
`STIMULI(5'h14, 5'h01, 5'h04, 32'h37890d6f, 1'h0)
`STIMULI(5'h18, 5'h0d, 5'h05, 32'he9d576d3, 1'h1)
`STIMULI(5'h08, 5'h05, 5'h06, 32'h7c99cff9, 1'h0)
`STIMULI(5'h03, 5'h10, 5'h07, 32'ha46c4848, 1'h1)
`STIMULI(5'h07, 5'h10, 5'h08, 32'h4506218a, 1'h0)
`STIMULI(5'h0e, 5'h0f, 5'h09, 32'h3058ef60, 1'h0)
`STIMULI(5'h12, 5'h14, 5'h0a, 32'hb955b672, 1'h0)
`STIMULI(5'h18, 5'h1e, 5'h0b, 32'hf40968e8, 1'h0)
`STIMULI(5'h0d, 5'h0b, 5'h0c, 32'h7c502bf8, 1'h1)
`STIMULI(5'h18, 5'h00, 5'h0d, 32'hd7e1c6af, 1'h0)
`STIMULI(5'h14, 5'h01, 5'h0e, 32'h50d909a1, 1'h1)
`STIMULI(5'h05, 5'h0b, 5'h0f, 32'h10c2c521, 1'h0)
`STIMULI(5'h0e, 5'h1c, 5'h10, 32'h1dd3013b, 1'h1)
`STIMULI(5'h00, 5'h02, 5'h11, 32'h0b636716, 1'h1)
`STIMULI(5'h0d, 5'h05, 5'h12, 32'hca91f895, 1'h0)
`STIMULI(5'h08, 5'h18, 5'h13, 32'h83a5a007, 1'h1)
`STIMULI(5'h17, 5'h0b, 5'h14, 32'h34243768, 1'h0)
`STIMULI(5'h12, 5'h03, 5'h15, 32'h9bcdf237, 1'h1)
`STIMULI(5'h11, 5'h14, 5'h16, 32'hc37a7886, 1'h1)
`STIMULI(5'h12, 5'h12, 5'h17, 32'hba460274, 1'h1)
`STIMULI(5'h08, 5'h04, 5'h18, 32'h66371fcc, 1'h0)
`STIMULI(5'h0c, 5'h14, 5'h19, 32'h41524b82, 1'h1)
`STIMULI(5'h05, 5'h01, 5'h1a, 32'hc7ac408f, 1'h1)
`STIMULI(5'h0b, 5'h16, 5'h1b, 32'h8ae2ac15, 1'h0)
`STIMULI(5'h15, 5'h1d, 5'h1c, 32'h1550d12a, 1'h0)
`STIMULI(5'h1b, 5'h0e, 5'h1d, 32'h23661746, 1'h1)
`STIMULI(5'h04, 5'h04, 5'h1e, 32'h49b4c193, 1'h1)
`STIMULI(5'h12, 5'h11, 5'h1f, 32'hb9492472, 1'h0)
`STIMULI(5'h03, 5'h0c, 5'h00, 32'h5abc1db5, 1'h0)
`STIMULI(5'h11, 5'h1e, 5'h01, 32'hcb87ba97, 1'h1)
`STIMULI(5'h16, 5'h14, 5'h02, 32'haba92e57, 1'h1)
`STIMULI(5'h13, 5'h09, 5'h03, 32'h8079ac00, 1'h0)
`STIMULI(5'h1e, 5'h0d, 5'h04, 32'h393d9b72, 1'h0)
`STIMULI(5'h1d, 5'h17, 5'h05, 32'h66c259cd, 1'h1)
`STIMULI(5'h0e, 5'h16, 5'h06, 32'h0dfa7f1b, 1'h0)
`STIMULI(5'h07, 5'h0d, 5'h07, 32'he50b48ca, 1'h0)
`STIMULI(5'h05, 5'h02, 5'h08, 32'h16479b2c, 1'h1)
`STIMULI(5'h03, 5'h1d, 5'h09, 32'hf9f1d4f3, 1'h1)
`STIMULI(5'h19, 5'h0c, 5'h0a, 32'h580965b0, 1'h0)
`STIMULI(5'h1a, 5'h02, 5'h0b, 32'h544fbfa8, 1'h0)
`STIMULI(5'h1c, 5'h1f, 5'h0c, 32'h4eee339d, 1'h1)
`STIMULI(5'h0c, 5'h00, 5'h0d, 32'hecc6d4d9, 1'h0)
`STIMULI(5'h01, 5'h0f, 5'h0e, 32'hae7a545c, 1'h0)
`STIMULI(5'h03, 5'h08, 5'h0f, 32'hd43790a8, 1'h1)
`STIMULI(5'h1d, 5'h18, 5'h10, 32'h7c9b37f9, 1'h1)
`STIMULI(5'h0b, 5'h1d, 5'h11, 32'h0f8abb1f, 1'h0)
`STIMULI(5'h0b, 5'h11, 5'h12, 32'h4b498396, 1'h1)
`STIMULI(5'h1f, 5'h0a, 5'h13, 32'hc7f6028f, 1'h0)
`STIMULI(5'h0d, 5'h05, 5'h14, 32'hbd823a7b, 1'h1)
`STIMULI(5'h1d, 5'h0a, 5'h15, 32'hffa3aaff, 1'h1)
`STIMULI(5'h1d, 5'h1d, 5'h16, 32'h6b9ee1d7, 1'h0)
`STIMULI(5'h0b, 5'h12, 5'h17, 32'h0d651b1a, 1'h1)
`STIMULI(5'h13, 5'h06, 5'h18, 32'h14d49329, 1'h1)
`STIMULI(5'h16, 5'h12, 5'h19, 32'h8ed88a1d, 1'h1)
`STIMULI(5'h12, 5'h17, 5'h1a, 32'hc762268e, 1'h0)
`STIMULI(5'h05, 5'h1e, 5'h1b, 32'hf7299aee, 1'h1)
`STIMULI(5'h07, 5'h04, 5'h1c, 32'hb6b5506d, 1'h1)
`STIMULI(5'h19, 5'h06, 5'h1d, 32'h9154fc22, 1'h1)
`STIMULI(5'h05, 5'h1b, 5'h1e, 32'hc68ec48d, 1'h0)
`STIMULI(5'h0c, 5'h0b, 5'h1f, 32'h679709cf, 1'h0)
`STIMULI(5'h18, 5'h03, 5'h00, 32'hd3ed4ca7, 1'h1)
`STIMULI(5'h0f, 5'h1b, 5'h01, 32'h366d676c, 1'h0)
`STIMULI(5'h0f, 5'h17, 5'h02, 32'h6847f1d0, 1'h0)
`STIMULI(5'h0e, 5'h05, 5'h03, 32'h1053a720, 1'h1)
`STIMULI(5'h14, 5'h04, 5'h04, 32'h395f1772, 1'h0)
`STIMULI(5'h13, 5'h03, 5'h05, 32'hd022e8a0, 1'h0)
`STIMULI(5'h1c, 5'h14, 5'h06, 32'h8fac9e1f, 1'h1)
`STIMULI(5'h04, 5'h0e, 5'h07, 32'h9abc7835, 1'h1)
`STIMULI(5'h19, 5'h04, 5'h08, 32'hd73b04ae, 1'h0)
`STIMULI(5'h0d, 5'h06, 5'h09, 32'had676c5a, 1'h1)
`STIMULI(5'h1c, 5'h01, 5'h0a, 32'h2a6b8354, 1'h0)
`STIMULI(5'h17, 5'h0b, 5'h0b, 32'h3d09457a, 1'h1)
`STIMULI(5'h19, 5'h1e, 5'h0c, 32'h03f32b07, 1'h1)
`STIMULI(5'h1b, 5'h05, 5'h0d, 32'h6b2191d6, 1'h1)
`STIMULI(5'h1b, 5'h08, 5'h0e, 32'h651711ca, 1'h1)
`STIMULI(5'h11, 5'h1c, 5'h0f, 32'h00308d00, 1'h0)
`STIMULI(5'h11, 5'h19, 5'h10, 32'h0eef5d1d, 1'h0)
`STIMULI(5'h11, 5'h0f, 5'h11, 32'hdff0bcbf, 1'h1)
`STIMULI(5'h1f, 5'h10, 5'h12, 32'he1397ac2, 1'h0)
`STIMULI(5'h18, 5'h17, 5'h13, 32'hba8b9475, 1'h1)
`STIMULI(5'h11, 5'h07, 5'h14, 32'h77012fee, 1'h0)
`STIMULI(5'h18, 5'h0f, 5'h15, 32'h86b1140d, 1'h1)
`STIMULI(5'h0b, 5'h14, 5'h16, 32'ha128b842, 1'h1)
`STIMULI(5'h1c, 5'h05, 5'h17, 32'h833a6206, 1'h0)
`STIMULI(5'h17, 5'h08, 5'h18, 32'hd897f4b1, 1'h0)
`STIMULI(5'h12, 5'h1e, 5'h19, 32'h0bbf7917, 1'h1)
`STIMULI(5'h0d, 5'h02, 5'h1a, 32'h1d9a7b3b, 1'h1)
`STIMULI(5'h1f, 5'h08, 5'h1b, 32'h2247b944, 1'h1)
`STIMULI(5'h12, 5'h00, 5'h1c, 32'h67b4c1cf, 1'h0)
`STIMULI(5'h17, 5'h19, 5'h1d, 32'h60fd93c1, 1'h0)
`STIMULI(5'h1f, 5'h16, 5'h1e, 32'hb8f83871, 1'h1)
`STIMULI(5'h06, 5'h0c, 5'h1f, 32'hc18d1c83, 1'h0)
`STIMULI(5'h10, 5'h0c, 5'h00, 32'h899e6a13, 1'h0)
`STIMULI(5'h1b, 5'h0e, 5'h01, 32'h7c95c1f9, 1'h1)
`STIMULI(5'h12, 5'h0d, 5'h02, 32'h84732208, 1'h1)
`STIMULI(5'h0d, 5'h0b, 5'h03, 32'he256d0c4, 1'h1)
`STIMULI(5'h0f, 5'h1d, 5'h04, 32'he25582c4, 1'h0)
`STIMULI(5'h03, 5'h1f, 5'h05, 32'ha67f2a4c, 1'h1)
`STIMULI(5'h0c, 5'h0e, 5'h06, 32'h0ad82f15, 1'h1)
`STIMULI(5'h19, 5'h16, 5'h07, 32'h5bc7d9b7, 1'h0)
`STIMULI(5'h00, 5'h13, 5'h08, 32'he9c860d3, 1'h0)
`STIMULI(5'h15, 5'h09, 5'h09, 32'hf8c1b2f1, 1'h0)
`STIMULI(5'h02, 5'h10, 5'h0a, 32'h9524102a, 1'h1)
`STIMULI(5'h15, 5'h17, 5'h0b, 32'he5fdfacb, 1'h1)
`STIMULI(5'h13, 5'h1a, 5'h0c, 32'hdcc714b9, 1'h1)
`STIMULI(5'h1c, 5'h12, 5'h0d, 32'h7679ffec, 1'h0)
`STIMULI(5'h00, 5'h0a, 5'h0e, 32'h1cd73d39, 1'h0)
`STIMULI(5'h0e, 5'h10, 5'h0f, 32'h75f5b9eb, 1'h0)
`STIMULI(5'h1d, 5'h18, 5'h10, 32'h9db7743b, 1'h1)
`STIMULI(5'h08, 5'h0b, 5'h11, 32'hdd9d70bb, 1'h1)
`STIMULI(5'h17, 5'h0e, 5'h12, 32'he009e4c0, 1'h1)
`STIMULI(5'h16, 5'h02, 5'h13, 32'h6e2e59dc, 1'h1)
`STIMULI(5'h08, 5'h03, 5'h14, 32'hd90912b2, 1'h0)
`STIMULI(5'h07, 5'h0a, 5'h15, 32'h177e2d2e, 1'h1)
`STIMULI(5'h01, 5'h04, 5'h16, 32'h4b400196, 1'h1)
`STIMULI(5'h01, 5'h19, 5'h17, 32'h680ddbd0, 1'h1)
`STIMULI(5'h1e, 5'h01, 5'h18, 32'h81694602, 1'h1)
`STIMULI(5'h06, 5'h04, 5'h19, 32'hec0f18d8, 1'h1)
`STIMULI(5'h04, 5'h1c, 5'h1a, 32'hacfd4059, 1'h1)
`STIMULI(5'h1a, 5'h1c, 5'h1b, 32'h1a050934, 1'h1)
`STIMULI(5'h15, 5'h00, 5'h1c, 32'h77b723ef, 1'h0)
`STIMULI(5'h07, 5'h16, 5'h1d, 32'h5be7d7b7, 1'h1)
`STIMULI(5'h1e, 5'h0c, 5'h1e, 32'he7191ace, 1'h0)
`STIMULI(5'h1a, 5'h0a, 5'h1f, 32'h9e73603c, 1'h0)
`STIMULI(5'h0b, 5'h1e, 5'h00, 32'hf2b778e5, 1'h0)
`STIMULI(5'h09, 5'h17, 5'h01, 32'hc508cc8a, 1'h1)
`STIMULI(5'h17, 5'h1c, 5'h02, 32'h11d2c523, 1'h1)
`STIMULI(5'h12, 5'h0a, 5'h03, 32'h1f4b2b3e, 1'h1)
`STIMULI(5'h02, 5'h05, 5'h04, 32'hfa88e0f5, 1'h1)
`STIMULI(5'h11, 5'h0d, 5'h05, 32'hb65f1c6c, 1'h1)
`STIMULI(5'h0f, 5'h0b, 5'h06, 32'hc4a52e89, 1'h1)
`STIMULI(5'h1b, 5'h00, 5'h07, 32'haa756854, 1'h1)
`STIMULI(5'h0f, 5'h03, 5'h08, 32'h0bd7ab17, 1'h1)
`STIMULI(5'h1c, 5'h1b, 5'h09, 32'h1608ab2c, 1'h1)
`STIMULI(5'h06, 5'h11, 5'h0a, 32'h78db0ff1, 1'h0)
`STIMULI(5'h14, 5'h1c, 5'h0b, 32'hb2f5e065, 1'h0)
`STIMULI(5'h13, 5'h00, 5'h0c, 32'hb6d1ec6d, 1'h0)
`STIMULI(5'h1f, 5'h00, 5'h0d, 32'hfe581afc, 1'h1)
`STIMULI(5'h0a, 5'h09, 5'h0e, 32'h39e2d773, 1'h0)
`STIMULI(5'h0e, 5'h05, 5'h0f, 32'h82cf1405, 1'h0)
`STIMULI(5'h0d, 5'h07, 5'h10, 32'hcddb7a9b, 1'h0)
`STIMULI(5'h1f, 5'h1f, 5'h11, 32'h7598d3eb, 1'h1)
`STIMULI(5'h15, 5'h0f, 5'h12, 32'h9762be2e, 1'h1)
`STIMULI(5'h17, 5'h07, 5'h13, 32'ha1a64a43, 1'h0)
`STIMULI(5'h11, 5'h01, 5'h14, 32'h7801e9f0, 1'h0)
`STIMULI(5'h09, 5'h0a, 5'h15, 32'he492f6c9, 1'h0)
`STIMULI(5'h1d, 5'h0f, 5'h16, 32'h8d0cb81a, 1'h1)
`STIMULI(5'h0d, 5'h17, 5'h17, 32'hf42782e8, 1'h1)
`STIMULI(5'h09, 5'h02, 5'h18, 32'h3b308b76, 1'h0)
`STIMULI(5'h0e, 5'h07, 5'h19, 32'hefcf68df, 1'h1)
`STIMULI(5'h02, 5'h16, 5'h1a, 32'hd43276a8, 1'h0)
`STIMULI(5'h12, 5'h1e, 5'h1b, 32'h18298730, 1'h1)
`STIMULI(5'h04, 5'h0b, 5'h1c, 32'hd22472a4, 1'h0)
`STIMULI(5'h16, 5'h01, 5'h1d, 32'h179bcd2f, 1'h0)
`STIMULI(5'h06, 5'h0f, 5'h1e, 32'hd3196ea6, 1'h0)
`STIMULI(5'h19, 5'h13, 5'h1f, 32'h4191d583, 1'h1)
`STIMULI(5'h00, 5'h06, 5'h00, 32'h622079c4, 1'h1)
`STIMULI(5'h03, 5'h0f, 5'h01, 32'h42ce8785, 1'h1)
`STIMULI(5'h0c, 5'h06, 5'h02, 32'h1e0ed53c, 1'h0)
`STIMULI(5'h14, 5'h0b, 5'h03, 32'h9bf8b437, 1'h1)
`STIMULI(5'h17, 5'h01, 5'h04, 32'h64612dc8, 1'h0)
`STIMULI(5'h15, 5'h09, 5'h05, 32'h184abd30, 1'h1)
`STIMULI(5'h11, 5'h0b, 5'h06, 32'h3e3b9d7c, 1'h0)
`STIMULI(5'h1c, 5'h00, 5'h07, 32'hf50d28ea, 1'h1)
`STIMULI(5'h15, 5'h00, 5'h08, 32'h5750e5ae, 1'h1)
`STIMULI(5'h1a, 5'h0c, 5'h09, 32'hcb445096, 1'h0)
`STIMULI(5'h1e, 5'h10, 5'h0a, 32'h32387b64, 1'h0)
`STIMULI(5'h09, 5'h09, 5'h0b, 32'h33b8f767, 1'h0)
`STIMULI(5'h1b, 5'h11, 5'h0c, 32'h0b7bb516, 1'h0)
`STIMULI(5'h0c, 5'h01, 5'h0d, 32'hbe43e87c, 1'h1)
`STIMULI(5'h08, 5'h12, 5'h0e, 32'hdc61e2b8, 1'h1)
`STIMULI(5'h1e, 5'h13, 5'h0f, 32'he004a0c0, 1'h0)
`STIMULI(5'h04, 5'h12, 5'h10, 32'h20437140, 1'h0)
`STIMULI(5'h1d, 5'h0f, 5'h11, 32'h20eae741, 1'h1)
`STIMULI(5'h13, 5'h0f, 5'h12, 32'h52ec09a5, 1'h0)
`STIMULI(5'h0f, 5'h1b, 5'h13, 32'hbfbb6c7f, 1'h1)
`STIMULI(5'h03, 5'h02, 5'h14, 32'h0453ad08, 1'h0)
`STIMULI(5'h13, 5'h17, 5'h15, 32'h6c776fd8, 1'h1)
`STIMULI(5'h14, 5'h10, 5'h16, 32'hc5b6de8b, 1'h1)
`STIMULI(5'h0c, 5'h1c, 5'h17, 32'h4bcf5b97, 1'h0)
`STIMULI(5'h12, 5'h14, 5'h18, 32'h8dd5bc1b, 1'h1)
`STIMULI(5'h00, 5'h00, 5'h19, 32'h630867c6, 1'h1)
`STIMULI(5'h07, 5'h1b, 5'h1a, 32'h6de21ddb, 1'h0)
`STIMULI(5'h18, 5'h07, 5'h1b, 32'h827d3404, 1'h0)
`STIMULI(5'h0b, 5'h01, 5'h1c, 32'hfe64b2fc, 1'h0)
`STIMULI(5'h08, 5'h19, 5'h1d, 32'hf5a170eb, 1'h0)
`STIMULI(5'h14, 5'h08, 5'h1e, 32'hbb213276, 1'h1)
`STIMULI(5'h0c, 5'h0b, 5'h1f, 32'h5a3079b4, 1'h1)
`STIMULI(5'h1f, 5'h0b, 5'h00, 32'h06c1670d, 1'h1)
`STIMULI(5'h0c, 5'h06, 5'h01, 32'h34eef369, 1'h1)
`STIMULI(5'h19, 5'h01, 5'h02, 32'hb2cf5665, 1'h1)
`STIMULI(5'h04, 5'h0e, 5'h03, 32'hd9276eb2, 1'h0)
`STIMULI(5'h12, 5'h0e, 5'h04, 32'h1e46693c, 1'h0)
`STIMULI(5'h01, 5'h06, 5'h05, 32'h30ca0f61, 1'h0)
`STIMULI(5'h12, 5'h02, 5'h06, 32'h34c37d69, 1'h0)
`STIMULI(5'h02, 5'h00, 5'h07, 32'h95d7182b, 1'h0)
`STIMULI(5'h16, 5'h0e, 5'h08, 32'h421c0f84, 1'h0)
`STIMULI(5'h02, 5'h03, 5'h09, 32'h6a7ca9d4, 1'h0)
`STIMULI(5'h17, 5'h13, 5'h0a, 32'h99e45833, 1'h1)
`STIMULI(5'h03, 5'h04, 5'h0b, 32'h240f3d48, 1'h1)
`STIMULI(5'h02, 5'h0a, 5'h0c, 32'hf02c6ee0, 1'h1)
`STIMULI(5'h02, 5'h1d, 5'h0d, 32'h3dc5677b, 1'h1)
`STIMULI(5'h02, 5'h0b, 5'h0e, 32'he07c5ec0, 1'h1)
`STIMULI(5'h04, 5'h0c, 5'h0f, 32'hb2de5c65, 1'h1)
`STIMULI(5'h1d, 5'h1a, 5'h10, 32'hf1d758e3, 1'h1)
`STIMULI(5'h00, 5'h17, 5'h11, 32'h649babc9, 1'h0)
`STIMULI(5'h06, 5'h01, 5'h12, 32'h5a4dc3b4, 1'h0)
`STIMULI(5'h09, 5'h0a, 5'h13, 32'hdf35bebe, 1'h0)
`STIMULI(5'h0d, 5'h00, 5'h14, 32'h4a666194, 1'h0)
`STIMULI(5'h14, 5'h10, 5'h15, 32'h79b399f3, 1'h0)
`STIMULI(5'h16, 5'h1a, 5'h16, 32'h90667620, 1'h0)
`STIMULI(5'h01, 5'h1f, 5'h17, 32'h7f4d65fe, 1'h1)
`STIMULI(5'h0a, 5'h16, 5'h18, 32'h5d40dfba, 1'h1)
`STIMULI(5'h07, 5'h03, 5'h19, 32'h1dc2173b, 1'h0)
`STIMULI(5'h0d, 5'h0d, 5'h1a, 32'hd0b432a1, 1'h1)
`STIMULI(5'h16, 5'h0a, 5'h1b, 32'heac812d5, 1'h0)
`STIMULI(5'h0e, 5'h19, 5'h1c, 32'h1fdfe53f, 1'h1)
`STIMULI(5'h19, 5'h13, 5'h1d, 32'h2380c747, 1'h1)
`STIMULI(5'h1b, 5'h17, 5'h1e, 32'h99586632, 1'h1)
`STIMULI(5'h15, 5'h10, 5'h1f, 32'h03974d07, 1'h0)
`STIMULI(5'h10, 5'h0c, 5'h00, 32'heb8244d7, 1'h0)
`STIMULI(5'h1f, 5'h05, 5'h01, 32'he6720ccc, 1'h0)
`STIMULI(5'h1c, 5'h1e, 5'h02, 32'hd5bc48ab, 1'h1)
`STIMULI(5'h0a, 5'h0a, 5'h03, 32'h039f5907, 1'h1)
`STIMULI(5'h0c, 5'h02, 5'h04, 32'h42a09785, 1'h0)
`STIMULI(5'h00, 5'h11, 5'h05, 32'hb0650e60, 1'h1)
`STIMULI(5'h0e, 5'h01, 5'h06, 32'ha164cc42, 1'h0)
`STIMULI(5'h0d, 5'h04, 5'h07, 32'hd31b3aa6, 1'h0)
`STIMULI(5'h10, 5'h0a, 5'h08, 32'h9e212a3c, 1'h0)
`STIMULI(5'h1a, 5'h1d, 5'h09, 32'hd1b9aea3, 1'h0)
`STIMULI(5'h16, 5'h19, 5'h0a, 32'h0486a709, 1'h0)
`STIMULI(5'h07, 5'h09, 5'h0b, 32'h6bc0b3d7, 1'h0)
`STIMULI(5'h19, 5'h1d, 5'h0c, 32'h164c172c, 1'h1)
`STIMULI(5'h1a, 5'h18, 5'h0d, 32'hd06492a0, 1'h0)
`STIMULI(5'h19, 5'h0f, 5'h0e, 32'hde5a4abc, 1'h0)
`STIMULI(5'h1d, 5'h19, 5'h0f, 32'h8ca44819, 1'h1)
`STIMULI(5'h0d, 5'h1a, 5'h10, 32'h7b7f2ff6, 1'h0)
`STIMULI(5'h00, 5'h0d, 5'h11, 32'hd1b31ca3, 1'h0)
`STIMULI(5'h18, 5'h12, 5'h12, 32'hf12feae2, 1'h1)
`STIMULI(5'h0b, 5'h18, 5'h13, 32'hc2dd4085, 1'h1)
`STIMULI(5'h14, 5'h0d, 5'h14, 32'h32a20765, 1'h1)
`STIMULI(5'h11, 5'h0d, 5'h15, 32'h22cf7145, 1'h0)
`STIMULI(5'h08, 5'h18, 5'h16, 32'hc4437e88, 1'h0)
`STIMULI(5'h08, 5'h11, 5'h17, 32'h8ae99c15, 1'h1)
`STIMULI(5'h1c, 5'h01, 5'h18, 32'he959f0d2, 1'h1)
`STIMULI(5'h09, 5'h1a, 5'h19, 32'h84047408, 1'h1)
`STIMULI(5'h05, 5'h04, 5'h1a, 32'hcf50b69e, 1'h1)
`STIMULI(5'h10, 5'h10, 5'h1b, 32'h0ed2211d, 1'h0)
`STIMULI(5'h0b, 5'h03, 5'h1c, 32'hf5fe04eb, 1'h1)
`STIMULI(5'h1c, 5'h1d, 5'h1d, 32'h9ac1ca35, 1'h1)
`STIMULI(5'h07, 5'h16, 5'h1e, 32'h23e70b47, 1'h1)
`STIMULI(5'h0c, 5'h16, 5'h1f, 32'hc50e508a, 1'h1)
`STIMULI(5'h12, 5'h1f, 5'h00, 32'hf74b14ee, 1'h0)
`STIMULI(5'h0e, 5'h0c, 5'h01, 32'hae5fd85c, 1'h1)
`STIMULI(5'h0d, 5'h04, 5'h02, 32'h887daa10, 1'h0)
`STIMULI(5'h07, 5'h10, 5'h03, 32'hf42872e8, 1'h0)
`STIMULI(5'h18, 5'h0a, 5'h04, 32'h07d7b30f, 1'h1)
`STIMULI(5'h12, 5'h0c, 5'h05, 32'h93a3c027, 1'h0)
`STIMULI(5'h16, 5'h0f, 5'h06, 32'hb9478c72, 1'h0)
`STIMULI(5'h13, 5'h06, 5'h07, 32'hdf218abe, 1'h1)
`STIMULI(5'h19, 5'h08, 5'h08, 32'h99483432, 1'h0)
`STIMULI(5'h05, 5'h11, 5'h09, 32'h6b0367d6, 1'h0)
`STIMULI(5'h18, 5'h16, 5'h0a, 32'h42c76585, 1'h0)
`STIMULI(5'h15, 5'h11, 5'h0b, 32'h1e95593d, 1'h0)
`STIMULI(5'h09, 5'h17, 5'h0c, 32'hcb42ae96, 1'h0)
`STIMULI(5'h03, 5'h0a, 5'h0d, 32'h95a9702b, 1'h0)
`STIMULI(5'h04, 5'h14, 5'h0e, 32'h2a23a754, 1'h1)
`STIMULI(5'h1f, 5'h1b, 5'h0f, 32'h6a9e65d5, 1'h1)
`STIMULI(5'h1f, 5'h03, 5'h10, 32'hd222f4a4, 1'h0)
`STIMULI(5'h0a, 5'h1c, 5'h11, 32'h0539410a, 1'h0)
`STIMULI(5'h0c, 5'h05, 5'h12, 32'h573a85ae, 1'h1)
`STIMULI(5'h10, 5'h00, 5'h13, 32'hd979f2b2, 1'h1)
`STIMULI(5'h18, 5'h12, 5'h14, 32'hc16e9a82, 1'h1)
`STIMULI(5'h08, 5'h1e, 5'h15, 32'hca52fa94, 1'h1)
`STIMULI(5'h08, 5'h0c, 5'h16, 32'h7475f7e8, 1'h1)
`STIMULI(5'h12, 5'h18, 5'h17, 32'h56ec05ad, 1'h1)
`STIMULI(5'h08, 5'h06, 5'h18, 32'hce08f49c, 1'h1)
`STIMULI(5'h03, 5'h08, 5'h19, 32'h85d7840b, 1'h0)
`STIMULI(5'h17, 5'h13, 5'h1a, 32'hb85fac70, 1'h1)
`STIMULI(5'h1f, 5'h1c, 5'h1b, 32'hd8635eb0, 1'h0)
`STIMULI(5'h16, 5'h06, 5'h1c, 32'hdc2714b8, 1'h0)
`STIMULI(5'h1d, 5'h1c, 5'h1d, 32'h20ec8141, 1'h0)
`STIMULI(5'h1d, 5'h15, 5'h1e, 32'hccf51e99, 1'h1)
`STIMULI(5'h03, 5'h0a, 5'h1f, 32'h91dd8423, 1'h1)
`STIMULI(5'h1c, 5'h12, 5'h00, 32'hed03d2da, 1'h0)
`STIMULI(5'h06, 5'h15, 5'h01, 32'hefc052df, 1'h1)
`STIMULI(5'h1b, 5'h13, 5'h02, 32'hc8bb7c91, 1'h1)
`STIMULI(5'h12, 5'h08, 5'h03, 32'h2f8abd5f, 1'h1)
`STIMULI(5'h02, 5'h0c, 5'h04, 32'hc053be80, 1'h0)
`STIMULI(5'h13, 5'h14, 5'h05, 32'h230e2146, 1'h0)
`STIMULI(5'h14, 5'h09, 5'h06, 32'hed93bcdb, 1'h0)
`STIMULI(5'h05, 5'h19, 5'h07, 32'hd8320ab0, 1'h0)
`STIMULI(5'h1e, 5'h15, 5'h08, 32'hbd792e7a, 1'h1)
`STIMULI(5'h1b, 5'h0f, 5'h09, 32'h2c61cf58, 1'h1)
`STIMULI(5'h12, 5'h1a, 5'h0a, 32'ha14e9242, 1'h1)
`STIMULI(5'h02, 5'h07, 5'h0b, 32'h7c552ff8, 1'h0)
`STIMULI(5'h12, 5'h1a, 5'h0c, 32'hf87838f0, 1'h1)
`STIMULI(5'h05, 5'h05, 5'h0d, 32'h791bfdf2, 1'h0)
`STIMULI(5'h13, 5'h06, 5'h0e, 32'hd40070a8, 1'h0)
`STIMULI(5'h16, 5'h0c, 5'h0f, 32'hb614b06c, 1'h0)
`STIMULI(5'h16, 5'h01, 5'h10, 32'he6aaaccd, 1'h0)
`STIMULI(5'h07, 5'h0a, 5'h11, 32'ha8361250, 1'h0)
`STIMULI(5'h1d, 5'h16, 5'h12, 32'hc8158e90, 1'h0)
`STIMULI(5'h0e, 5'h18, 5'h13, 32'h3dd3d57b, 1'h0)
`STIMULI(5'h0f, 5'h0f, 5'h14, 32'h17341f2e, 1'h1)
`STIMULI(5'h0e, 5'h09, 5'h15, 32'h1ec6353d, 1'h0)
`STIMULI(5'h0d, 5'h12, 5'h16, 32'hf025dee0, 1'h0)
`STIMULI(5'h0d, 5'h13, 5'h17, 32'hb79c9c6f, 1'h1)
`STIMULI(5'h07, 5'h0c, 5'h18, 32'h0335e706, 1'h1)
`STIMULI(5'h09, 5'h06, 5'h19, 32'h9f43423e, 1'h1)
`STIMULI(5'h05, 5'h04, 5'h1a, 32'h568913ad, 1'h1)
`STIMULI(5'h16, 5'h08, 5'h1b, 32'h5d43cdba, 1'h1)
`STIMULI(5'h1b, 5'h00, 5'h1c, 32'hc9c31693, 1'h0)
`STIMULI(5'h00, 5'h0d, 5'h1d, 32'h4788e78f, 1'h0)
`STIMULI(5'h18, 5'h1c, 5'h1e, 32'hc2aaa085, 1'h0)
`STIMULI(5'h04, 5'h12, 5'h1f, 32'hc94ce892, 1'h0)
`STIMULI(5'h1f, 5'h0c, 5'h00, 32'h6b9481d7, 1'h1)
`STIMULI(5'h07, 5'h0f, 5'h01, 32'h199b7f33, 1'h1)
`STIMULI(5'h0c, 5'h03, 5'h02, 32'h901dbc20, 1'h0)
`STIMULI(5'h1c, 5'h12, 5'h03, 32'he68e36cd, 1'h0)
`STIMULI(5'h0a, 5'h04, 5'h04, 32'hda7cbcb4, 1'h1)
`STIMULI(5'h13, 5'h1c, 5'h05, 32'hf32c32e6, 1'h1)
`STIMULI(5'h0a, 5'h07, 5'h06, 32'heb715cd6, 1'h1)
`STIMULI(5'h09, 5'h09, 5'h07, 32'hc894ba91, 1'h1)
`STIMULI(5'h05, 5'h15, 5'h08, 32'hf09c1ae1, 1'h1)
`STIMULI(5'h0d, 5'h1b, 5'h09, 32'h97dce42f, 1'h0)
`STIMULI(5'h12, 5'h09, 5'h0a, 32'he8c42ed1, 1'h0)
`STIMULI(5'h1d, 5'h14, 5'h0b, 32'hf0c834e1, 1'h0)
`STIMULI(5'h0c, 5'h02, 5'h0c, 32'h2354b146, 1'h1)
`STIMULI(5'h00, 5'h12, 5'h0d, 32'h32443b64, 1'h0)
`STIMULI(5'h0f, 5'h0b, 5'h0e, 32'ha818ac50, 1'h1)
`STIMULI(5'h09, 5'h1b, 5'h0f, 32'h444f2d88, 1'h0)
`STIMULI(5'h0e, 5'h15, 5'h10, 32'h85fe520b, 1'h0)
`STIMULI(5'h14, 5'h12, 5'h11, 32'h6fb197df, 1'h0)
`STIMULI(5'h1e, 5'h19, 5'h12, 32'h7b6909f6, 1'h0)
`STIMULI(5'h0f, 5'h0a, 5'h13, 32'hb6b2e66d, 1'h0)
`STIMULI(5'h08, 5'h1f, 5'h14, 32'h705a95e0, 1'h1)
`STIMULI(5'h13, 5'h0f, 5'h15, 32'h1ab11d35, 1'h0)
`STIMULI(5'h04, 5'h1c, 5'h16, 32'hc27b3484, 1'h1)
`STIMULI(5'h1a, 5'h19, 5'h17, 32'h6d4365da, 1'h1)
`STIMULI(5'h0d, 5'h14, 5'h18, 32'hdcc8c8b9, 1'h0)
`STIMULI(5'h09, 5'h09, 5'h19, 32'hd84fb2b0, 1'h1)
`STIMULI(5'h08, 5'h19, 5'h1a, 32'hf074e8e0, 1'h1)
`STIMULI(5'h1f, 5'h05, 5'h1b, 32'hdf3b6abe, 1'h0)
`STIMULI(5'h1f, 5'h0a, 5'h1c, 32'h523a07a4, 1'h1)
`STIMULI(5'h01, 5'h06, 5'h1d, 32'h6c1efbd8, 1'h0)
`STIMULI(5'h0d, 5'h0d, 5'h1e, 32'hef2f94de, 1'h1)
`STIMULI(5'h10, 5'h0b, 5'h1f, 32'h36a47f6d, 1'h1)
`STIMULI(5'h01, 5'h0a, 5'h00, 32'hede51edb, 1'h0)
`STIMULI(5'h0e, 5'h03, 5'h01, 32'ha6f95a4d, 1'h0)
`STIMULI(5'h00, 5'h03, 5'h02, 32'hd44c6ea8, 1'h1)
`STIMULI(5'h0e, 5'h05, 5'h03, 32'hf5fae0eb, 1'h1)
`STIMULI(5'h0d, 5'h08, 5'h04, 32'he0baa8c1, 1'h0)
`STIMULI(5'h1c, 5'h0e, 5'h05, 32'he485f2c9, 1'h0)
`STIMULI(5'h13, 5'h18, 5'h06, 32'h9c086a38, 1'h0)
`STIMULI(5'h1f, 5'h19, 5'h07, 32'ha6919a4d, 1'h0)
`STIMULI(5'h0b, 5'h03, 5'h08, 32'h7498f5e9, 1'h1)
`STIMULI(5'h03, 5'h16, 5'h09, 32'hbb7cac76, 1'h1)
`STIMULI(5'h1c, 5'h01, 5'h0a, 32'h5dd03dbb, 1'h1)
`STIMULI(5'h0c, 5'h14, 5'h0b, 32'h13b66b27, 1'h0)
`STIMULI(5'h09, 5'h02, 5'h0c, 32'h6d4019da, 1'h0)
`STIMULI(5'h0b, 5'h13, 5'h0d, 32'h44aa2789, 1'h1)
`STIMULI(5'h18, 5'h1f, 5'h0e, 32'h2e94595d, 1'h1)
`STIMULI(5'h14, 5'h12, 5'h0f, 32'h5695dbad, 1'h1)
`STIMULI(5'h1b, 5'h1b, 5'h10, 32'h5905e9b2, 1'h1)
`STIMULI(5'h09, 5'h0a, 5'h11, 32'h1cb3c939, 1'h0)
`STIMULI(5'h1b, 5'h19, 5'h12, 32'ha4dcf249, 1'h0)
`STIMULI(5'h19, 5'h1b, 5'h13, 32'hb6df286d, 1'h1)
`STIMULI(5'h09, 5'h13, 5'h14, 32'h2549f94a, 1'h1)
`STIMULI(5'h1a, 5'h08, 5'h15, 32'h049bb709, 1'h0)
`STIMULI(5'h13, 5'h15, 5'h16, 32'hb29dfc65, 1'h0)
`STIMULI(5'h17, 5'h19, 5'h17, 32'h24285d48, 1'h1)
`STIMULI(5'h02, 5'h16, 5'h18, 32'h0aa99d15, 1'h0)
`STIMULI(5'h06, 5'h19, 5'h19, 32'hc504d08a, 1'h1)
`STIMULI(5'h10, 5'h0a, 5'h1a, 32'h48cb2f91, 1'h0)
`STIMULI(5'h1c, 5'h1e, 5'h1b, 32'hcc123898, 1'h1)
`STIMULI(5'h1f, 5'h13, 5'h1c, 32'ha4f3e649, 1'h1)
`STIMULI(5'h13, 5'h16, 5'h1d, 32'hb836c070, 1'h0)
`STIMULI(5'h08, 5'h01, 5'h1e, 32'hf8abf8f1, 1'h0)
`STIMULI(5'h1f, 5'h09, 5'h1f, 32'h112c4322, 1'h0)
`STIMULI(5'h03, 5'h03, 5'h00, 32'hcaddae95, 1'h0)
`STIMULI(5'h0d, 5'h12, 5'h01, 32'h1ee1e53d, 1'h0)
`STIMULI(5'h0e, 5'h1d, 5'h02, 32'h86ef900d, 1'h1)
`STIMULI(5'h07, 5'h13, 5'h03, 32'he698bccd, 1'h0)
`STIMULI(5'h1c, 5'h05, 5'h04, 32'h797585f2, 1'h1)
`STIMULI(5'h11, 5'h10, 5'h05, 32'h23a36547, 1'h0)
`STIMULI(5'h00, 5'h02, 5'h06, 32'h2480eb49, 1'h0)
`STIMULI(5'h1e, 5'h03, 5'h07, 32'h5470aba8, 1'h0)
`STIMULI(5'h07, 5'h15, 5'h08, 32'he757bece, 1'h1)
`STIMULI(5'h1f, 5'h15, 5'h09, 32'h31492362, 1'h0)
`STIMULI(5'h0d, 5'h19, 5'h0a, 32'hc11aba82, 1'h0)
`STIMULI(5'h0e, 5'h1e, 5'h0b, 32'ha8e7d251, 1'h1)
`STIMULI(5'h11, 5'h05, 5'h0c, 32'h93a27027, 1'h0)
`STIMULI(5'h17, 5'h02, 5'h0d, 32'hffd5c4ff, 1'h1)
`STIMULI(5'h05, 5'h17, 5'h0e, 32'hab9b7457, 1'h1)
`STIMULI(5'h0c, 5'h13, 5'h0f, 32'h9a30b634, 1'h1)
`STIMULI(5'h08, 5'h03, 5'h10, 32'he4a96ec9, 1'h1)
`STIMULI(5'h14, 5'h1e, 5'h11, 32'h7c44adf8, 1'h1)
`STIMULI(5'h16, 5'h1b, 5'h12, 32'h74194de8, 1'h0)
`STIMULI(5'h08, 5'h07, 5'h13, 32'h5d209bba, 1'h1)
`STIMULI(5'h11, 5'h13, 5'h14, 32'haa6a4c54, 1'h1)
`STIMULI(5'h03, 5'h02, 5'h15, 32'h6f0dffde, 1'h0)
`STIMULI(5'h19, 5'h00, 5'h16, 32'hc3b63487, 1'h0)
`STIMULI(5'h15, 5'h1a, 5'h17, 32'h749385e9, 1'h1)
`STIMULI(5'h07, 5'h02, 5'h18, 32'h98c05e31, 1'h0)
`STIMULI(5'h1f, 5'h1b, 5'h19, 32'h856aa00a, 1'h1)
`STIMULI(5'h07, 5'h0b, 5'h1a, 32'h9e33e23c, 1'h1)
`STIMULI(5'h08, 5'h14, 5'h1b, 32'hbd90367b, 1'h1)
`STIMULI(5'h0f, 5'h01, 5'h1c, 32'h8d58b81a, 1'h1)
`STIMULI(5'h03, 5'h01, 5'h1d, 32'h21583542, 1'h1)
`STIMULI(5'h0c, 5'h08, 5'h1e, 32'h4147cd82, 1'h0)
`STIMULI(5'h04, 5'h1a, 5'h1f, 32'hfc2c36f8, 1'h1)
`STIMULI(5'h1c, 5'h05, 5'h00, 32'h35662d6a, 1'h0)
`STIMULI(5'h0f, 5'h13, 5'h01, 32'h145d2128, 1'h1)
`STIMULI(5'h05, 5'h0e, 5'h02, 32'h95af222b, 1'h0)
`STIMULI(5'h00, 5'h03, 5'h03, 32'hed2fc6da, 1'h1)
`STIMULI(5'h02, 5'h01, 5'h04, 32'h671551ce, 1'h1)
`STIMULI(5'h0b, 5'h1c, 5'h05, 32'h290c8752, 1'h0)
`STIMULI(5'h1c, 5'h05, 5'h06, 32'he602dacc, 1'h0)
`STIMULI(5'h16, 5'h1b, 5'h07, 32'ha079ea40, 1'h0)
`STIMULI(5'h05, 5'h17, 5'h08, 32'h42c07b85, 1'h0)
`STIMULI(5'h19, 5'h08, 5'h09, 32'h1f4a4b3e, 1'h1)
`STIMULI(5'h1b, 5'h1d, 5'h0a, 32'h4f4ba99e, 1'h1)
`STIMULI(5'h19, 5'h00, 5'h0b, 32'ha0246840, 1'h0)
`STIMULI(5'h04, 5'h0f, 5'h0c, 32'hefe3badf, 1'h0)
`STIMULI(5'h0c, 5'h10, 5'h0d, 32'h7f4f11fe, 1'h1)
`STIMULI(5'h08, 5'h1f, 5'h0e, 32'h1f56013e, 1'h1)
`STIMULI(5'h00, 5'h15, 5'h0f, 32'h2867c350, 1'h1)
`STIMULI(5'h18, 5'h19, 5'h10, 32'h89d0e613, 1'h1)
`STIMULI(5'h1d, 5'h12, 5'h11, 32'h676c3fce, 1'h1)
`STIMULI(5'h0a, 5'h1b, 5'h12, 32'h14c61529, 1'h0)
`STIMULI(5'h0f, 5'h02, 5'h13, 32'h743f3de8, 1'h0)
`STIMULI(5'h16, 5'h02, 5'h14, 32'h90239220, 1'h0)
`STIMULI(5'h03, 5'h05, 5'h15, 32'h388ff971, 1'h0)
`STIMULI(5'h0b, 5'h18, 5'h16, 32'h34ebdd69, 1'h1)
`STIMULI(5'h00, 5'h1c, 5'h17, 32'he2ccdcc5, 1'h0)
`STIMULI(5'h17, 5'h02, 5'h18, 32'heef510dd, 1'h0)
`STIMULI(5'h07, 5'h08, 5'h19, 32'hc589208b, 1'h1)
`STIMULI(5'h0f, 5'h05, 5'h1a, 32'hab570856, 1'h0)
`STIMULI(5'h15, 5'h03, 5'h1b, 32'h797d65f2, 1'h1)
`STIMULI(5'h1b, 5'h15, 5'h1c, 32'h72d079e5, 1'h0)
`STIMULI(5'h14, 5'h04, 5'h1d, 32'h690b5bd2, 1'h0)
`STIMULI(5'h16, 5'h0b, 5'h1e, 32'he72b10ce, 1'h1)
`STIMULI(5'h08, 5'h03, 5'h1f, 32'h06ec5b0d, 1'h0)
`STIMULI(5'h1b, 5'h17, 5'h00, 32'h3c669b78, 1'h0)
`STIMULI(5'h16, 5'h19, 5'h01, 32'h26730b4c, 1'h0)
`STIMULI(5'h0c, 5'h10, 5'h02, 32'hea3324d4, 1'h0)
`STIMULI(5'h0a, 5'h15, 5'h03, 32'hea8800d5, 1'h1)
`STIMULI(5'h01, 5'h19, 5'h04, 32'h88020e10, 1'h0)
`STIMULI(5'h1c, 5'h06, 5'h05, 32'hb9495672, 1'h1)
`STIMULI(5'h08, 5'h16, 5'h06, 32'h7db63bfb, 1'h1)
`STIMULI(5'h0d, 5'h0c, 5'h07, 32'h44f55b89, 1'h0)
`STIMULI(5'h0b, 5'h0c, 5'h08, 32'hdcbb24b9, 1'h0)
`STIMULI(5'h02, 5'h14, 5'h09, 32'h3788216f, 1'h1)
`STIMULI(5'h12, 5'h15, 5'h0a, 32'hc10b0682, 1'h0)
`STIMULI(5'h1a, 5'h00, 5'h0b, 32'h15342f2a, 1'h1)
`STIMULI(5'h1b, 5'h1b, 5'h0c, 32'h776bf3ee, 1'h1)
`STIMULI(5'h08, 5'h07, 5'h0d, 32'haa9e0e55, 1'h1)
`STIMULI(5'h07, 5'h1d, 5'h0e, 32'h45ebfb8b, 1'h1)
`STIMULI(5'h14, 5'h0b, 5'h0f, 32'h8682fe0d, 1'h0)
`STIMULI(5'h08, 5'h1f, 5'h10, 32'h85644c0a, 1'h1)
`STIMULI(5'h02, 5'h04, 5'h11, 32'hc3328286, 1'h0)
`STIMULI(5'h0b, 5'h0b, 5'h12, 32'hae8b4e5d, 1'h0)
`STIMULI(5'h1c, 5'h19, 5'h13, 32'h73030fe6, 1'h1)
`STIMULI(5'h06, 5'h18, 5'h14, 32'h82ddc605, 1'h1)
`STIMULI(5'h07, 5'h11, 5'h15, 32'h8ba9a017, 1'h1)
`STIMULI(5'h18, 5'h0f, 5'h16, 32'h8166f402, 1'h0)
`STIMULI(5'h1b, 5'h15, 5'h17, 32'hdf1c64be, 1'h1)
`STIMULI(5'h03, 5'h15, 5'h18, 32'hd12fb4a2, 1'h1)
`STIMULI(5'h0b, 5'h13, 5'h19, 32'hbd684e7a, 1'h1)
`STIMULI(5'h1f, 5'h1a, 5'h1a, 32'ha6dc9e4d, 1'h1)
`STIMULI(5'h0d, 5'h1b, 5'h1b, 32'hf1a1c2e3, 1'h1)
`STIMULI(5'h09, 5'h06, 5'h1c, 32'h58c329b1, 1'h1)
`STIMULI(5'h02, 5'h16, 5'h1d, 32'h1cd82f39, 1'h0)
`STIMULI(5'h1a, 5'h0b, 5'h1e, 32'hc47dc288, 1'h1)
`STIMULI(5'h0b, 5'h01, 5'h1f, 32'hacb4ae59, 1'h0)
`STIMULI(5'h08, 5'h17, 5'h00, 32'hcac6fa95, 1'h0)
`STIMULI(5'h1d, 5'h0b, 5'h01, 32'h002ba700, 1'h0)
`STIMULI(5'h02, 5'h12, 5'h02, 32'h6a2397d4, 1'h1)
`STIMULI(5'h0c, 5'h01, 5'h03, 32'h6b696bd6, 1'h0)
`STIMULI(5'h15, 5'h01, 5'h04, 32'hd6a3baad, 1'h1)
`STIMULI(5'h0e, 5'h1a, 5'h05, 32'he4e1d8c9, 1'h0)
`STIMULI(5'h1f, 5'h06, 5'h06, 32'hc4c30a89, 1'h1)
`STIMULI(5'h04, 5'h19, 5'h07, 32'he82afad0, 1'h0)
`STIMULI(5'h16, 5'h12, 5'h08, 32'h672fbfce, 1'h0)
`STIMULI(5'h03, 5'h18, 5'h09, 32'hb80aa870, 1'h0)
`STIMULI(5'h18, 5'h1d, 5'h0a, 32'h4b00d396, 1'h0)
`STIMULI(5'h19, 5'h1b, 5'h0b, 32'h4fdf259f, 1'h1)
`STIMULI(5'h07, 5'h1c, 5'h0c, 32'hbba31a77, 1'h0)
`STIMULI(5'h04, 5'h07, 5'h0d, 32'h354abd6a, 1'h0)
`STIMULI(5'h03, 5'h0e, 5'h0e, 32'h9785662f, 1'h1)
`STIMULI(5'h06, 5'h1e, 5'h0f, 32'ha5ca6a4b, 1'h0)
`STIMULI(5'h0b, 5'h0f, 5'h10, 32'hf04ba2e0, 1'h1)
`STIMULI(5'h19, 5'h07, 5'h11, 32'h809f7601, 1'h0)
`STIMULI(5'h04, 5'h18, 5'h12, 32'h6510f9ca, 1'h0)
`STIMULI(5'h13, 5'h0e, 5'h13, 32'h7c3411f8, 1'h1)
`STIMULI(5'h0a, 5'h07, 5'h14, 32'h4b00eb96, 1'h1)
`STIMULI(5'h16, 5'h1e, 5'h15, 32'hdee2fabd, 1'h0)
`STIMULI(5'h05, 5'h11, 5'h16, 32'h604f7bc0, 1'h0)
`STIMULI(5'h02, 5'h14, 5'h17, 32'hc5ca1c8b, 1'h1)
`STIMULI(5'h14, 5'h13, 5'h18, 32'h5f5847be, 1'h1)
`STIMULI(5'h11, 5'h06, 5'h19, 32'h31102f62, 1'h0)
`STIMULI(5'h0a, 5'h03, 5'h1a, 32'h436ca586, 1'h1)
`STIMULI(5'h13, 5'h08, 5'h1b, 32'h43c55187, 1'h1)
`STIMULI(5'h15, 5'h02, 5'h1c, 32'hde98cabd, 1'h1)
`STIMULI(5'h00, 5'h04, 5'h1d, 32'h9646b42c, 1'h1)
`STIMULI(5'h04, 5'h01, 5'h1e, 32'h6f67e7de, 1'h0)
`STIMULI(5'h08, 5'h08, 5'h1f, 32'hd4cd32a9, 1'h1)
`STIMULI(5'h03, 5'h1c, 5'h00, 32'ha76f484e, 1'h0)
`STIMULI(5'h18, 5'h0a, 5'h01, 32'h588ef1b1, 1'h0)
`STIMULI(5'h1e, 5'h1b, 5'h02, 32'hf72876ee, 1'h1)
`STIMULI(5'h07, 5'h17, 5'h03, 32'ha89c0451, 1'h1)
`STIMULI(5'h0f, 5'h09, 5'h04, 32'h696257d2, 1'h0)
`STIMULI(5'h02, 5'h1b, 5'h05, 32'h085e0910, 1'h1)
`STIMULI(5'h13, 5'h1a, 5'h06, 32'hd05148a0, 1'h1)
`STIMULI(5'h11, 5'h1c, 5'h07, 32'h1c62cb38, 1'h0)
`STIMULI(5'h1d, 5'h1d, 5'h08, 32'hf0064ae0, 1'h1)
`STIMULI(5'h1d, 5'h0c, 5'h09, 32'h6ad9e1d5, 1'h1)
`STIMULI(5'h0a, 5'h0c, 5'h0a, 32'h9dd5103b, 1'h1)
`STIMULI(5'h14, 5'h09, 5'h0b, 32'hc3ed4a87, 1'h0)
`STIMULI(5'h10, 5'h1e, 5'h0c, 32'he9f134d3, 1'h1)
`STIMULI(5'h11, 5'h0c, 5'h0d, 32'h9edd183d, 1'h0)
`STIMULI(5'h13, 5'h05, 5'h0e, 32'h484a4390, 1'h1)
`STIMULI(5'h0a, 5'h0e, 5'h0f, 32'he38606c7, 1'h0)
`STIMULI(5'h0c, 5'h1b, 5'h10, 32'hbf6eea7e, 1'h0)
`STIMULI(5'h12, 5'h08, 5'h11, 32'h9cbb1839, 1'h0)
`STIMULI(5'h17, 5'h06, 5'h12, 32'h57ff13af, 1'h0)
`STIMULI(5'h10, 5'h1f, 5'h13, 32'h5e9a43bd, 1'h0)
`STIMULI(5'h1e, 5'h18, 5'h14, 32'hccf50099, 1'h0)
`STIMULI(5'h0e, 5'h1a, 5'h15, 32'hf4c404e9, 1'h0)
`STIMULI(5'h11, 5'h1f, 5'h16, 32'hc4cd7289, 1'h0)
`STIMULI(5'h08, 5'h01, 5'h17, 32'hdf1e04be, 1'h0)
`STIMULI(5'h0c, 5'h0d, 5'h18, 32'h1556c92a, 1'h1)
`STIMULI(5'h15, 5'h05, 5'h19, 32'h7088bde1, 1'h1)
`STIMULI(5'h17, 5'h13, 5'h1a, 32'hafaf1a5f, 1'h1)
`STIMULI(5'h00, 5'h0a, 5'h1b, 32'hb9b00e73, 1'h0)
`STIMULI(5'h13, 5'h12, 5'h1c, 32'h3fb95b7f, 1'h0)
`STIMULI(5'h1c, 5'h14, 5'h1d, 32'hfadee8f5, 1'h0)
`STIMULI(5'h18, 5'h1d, 5'h1e, 32'h3a117b74, 1'h1)
`STIMULI(5'h10, 5'h07, 5'h1f, 32'hd27de6a4, 1'h1)
`STIMULI(5'h03, 5'h13, 5'h00, 32'h754787ea, 1'h0)
`STIMULI(5'h11, 5'h0f, 5'h01, 32'hf2a4ece5, 1'h1)
`STIMULI(5'h0f, 5'h0d, 5'h02, 32'h6ee9c9dd, 1'h1)
`STIMULI(5'h13, 5'h1f, 5'h03, 32'h86e7ce0d, 1'h1)
`STIMULI(5'h1b, 5'h14, 5'h04, 32'h72a5e5e5, 1'h0)
`STIMULI(5'h12, 5'h05, 5'h05, 32'hcc45ea98, 1'h0)
`STIMULI(5'h0d, 5'h12, 5'h06, 32'hf188f8e3, 1'h1)
`STIMULI(5'h03, 5'h0a, 5'h07, 32'h5fe4cbbf, 1'h1)
`STIMULI(5'h0d, 5'h18, 5'h08, 32'he126c4c2, 1'h0)
`STIMULI(5'h08, 5'h1c, 5'h09, 32'ha5fdc64b, 1'h0)
`STIMULI(5'h1c, 5'h0f, 5'h0a, 32'he62fbecc, 1'h0)
`STIMULI(5'h01, 5'h17, 5'h0b, 32'h1126a122, 1'h0)
`STIMULI(5'h16, 5'h03, 5'h0c, 32'hcbbe3c97, 1'h1)
`STIMULI(5'h14, 5'h06, 5'h0d, 32'h32dd2765, 1'h0)
`STIMULI(5'h09, 5'h11, 5'h0e, 32'h48628f90, 1'h1)
`STIMULI(5'h0f, 5'h15, 5'h0f, 32'h08fdd311, 1'h1)
`STIMULI(5'h0e, 5'h0e, 5'h10, 32'hc3b62087, 1'h0)
`STIMULI(5'h14, 5'h0c, 5'h11, 32'h208d6d41, 1'h1)
`STIMULI(5'h00, 5'h10, 5'h12, 32'ha2fd9c45, 1'h0)
`STIMULI(5'h08, 5'h00, 5'h13, 32'h94fda429, 1'h1)
`STIMULI(5'h1a, 5'h0d, 5'h14, 32'h09220512, 1'h1)
`STIMULI(5'h04, 5'h0e, 5'h15, 32'hdbd4bcb7, 1'h0)
`STIMULI(5'h12, 5'h16, 5'h16, 32'hde08dabc, 1'h1)
`STIMULI(5'h19, 5'h1a, 5'h17, 32'h5f601dbe, 1'h1)
`STIMULI(5'h05, 5'h0b, 5'h18, 32'hcb133c96, 1'h1)
`STIMULI(5'h0c, 5'h09, 5'h19, 32'h57d9fdaf, 1'h1)
`STIMULI(5'h09, 5'h13, 5'h1a, 32'h964c002c, 1'h0)
`STIMULI(5'h08, 5'h1d, 5'h1b, 32'hc929fc92, 1'h1)
`STIMULI(5'h10, 5'h14, 5'h1c, 32'h538cdba7, 1'h0)
`STIMULI(5'h18, 5'h03, 5'h1d, 32'h3c28cf78, 1'h1)
`STIMULI(5'h12, 5'h09, 5'h1e, 32'h32a27f65, 1'h0)
`STIMULI(5'h0b, 5'h02, 5'h1f, 32'h650ecbca, 1'h0)
`STIMULI(5'h18, 5'h03, 5'h00, 32'hb337b666, 1'h0)
`STIMULI(5'h0b, 5'h0a, 5'h01, 32'h9d75983a, 1'h0)
`STIMULI(5'h1c, 5'h1d, 5'h02, 32'hab0f8a56, 1'h1)
`STIMULI(5'h01, 5'h1a, 5'h03, 32'h9714c82e, 1'h0)
`STIMULI(5'h1b, 5'h01, 5'h04, 32'h40d66181, 1'h1)
`STIMULI(5'h11, 5'h0b, 5'h05, 32'h25217b4a, 1'h0)
`STIMULI(5'h10, 5'h04, 5'h06, 32'hb592186b, 1'h0)
`STIMULI(5'h02, 5'h0d, 5'h07, 32'h1cf8fb39, 1'h1)
`STIMULI(5'h0b, 5'h09, 5'h08, 32'h00792f00, 1'h1)
`STIMULI(5'h16, 5'h11, 5'h09, 32'h4b7e5f96, 1'h1)
`STIMULI(5'h1c, 5'h0c, 5'h0a, 32'hccb8dc99, 1'h1)
`STIMULI(5'h0e, 5'h0b, 5'h0b, 32'h03532706, 1'h0)
`STIMULI(5'h13, 5'h08, 5'h0c, 32'hc672348c, 1'h1)
`STIMULI(5'h0f, 5'h1f, 5'h0d, 32'h08d2e311, 1'h1)
`STIMULI(5'h0c, 5'h15, 5'h0e, 32'h43f64b87, 1'h1)
`STIMULI(5'h19, 5'h03, 5'h0f, 32'h4b79cf96, 1'h0)
`STIMULI(5'h0f, 5'h0b, 5'h10, 32'haa094654, 1'h0)
`STIMULI(5'h1d, 5'h0f, 5'h11, 32'h211e6f42, 1'h1)
`STIMULI(5'h11, 5'h0b, 5'h12, 32'h5db495bb, 1'h1)
`STIMULI(5'h06, 5'h1b, 5'h13, 32'h4626378c, 1'h1)
`STIMULI(5'h0c, 5'h1e, 5'h14, 32'h1beff937, 1'h0)
`STIMULI(5'h06, 5'h19, 5'h15, 32'hee9d26dd, 1'h1)
`STIMULI(5'h16, 5'h07, 5'h16, 32'h1729b32e, 1'h1)
`STIMULI(5'h17, 5'h17, 5'h17, 32'h66d865cd, 1'h0)
`STIMULI(5'h0f, 5'h0d, 5'h18, 32'hb4759e68, 1'h0)
`STIMULI(5'h02, 5'h06, 5'h19, 32'h4f0beb9e, 1'h1)
`STIMULI(5'h18, 5'h05, 5'h1a, 32'h1deb553b, 1'h0)
`STIMULI(5'h14, 5'h11, 5'h1b, 32'h13fb1b27, 1'h0)
`STIMULI(5'h10, 5'h01, 5'h1c, 32'h8d7b4a1a, 1'h1)
`STIMULI(5'h10, 5'h07, 5'h1d, 32'h17ac652f, 1'h1)
`STIMULI(5'h06, 5'h05, 5'h1e, 32'h2342f346, 1'h0)
`STIMULI(5'h1c, 5'h16, 5'h1f, 32'hb7c7de6f, 1'h0)
`STIMULI(5'h09, 5'h0a, 5'h00, 32'hbc27d478, 1'h1)
`STIMULI(5'h01, 5'h03, 5'h01, 32'h3408f368, 1'h0)
`STIMULI(5'h05, 5'h1d, 5'h02, 32'h8141bc02, 1'h0)
`STIMULI(5'h18, 5'h00, 5'h03, 32'h15eaf32b, 1'h0)
`STIMULI(5'h09, 5'h03, 5'h04, 32'h3e5bcd7c, 1'h1)
`STIMULI(5'h08, 5'h19, 5'h05, 32'h5378bda6, 1'h1)
`STIMULI(5'h16, 5'h1f, 5'h06, 32'he594a8cb, 1'h1)
`STIMULI(5'h0e, 5'h08, 5'h07, 32'ha9e75a53, 1'h1)
`STIMULI(5'h15, 5'h0b, 5'h08, 32'h6fe58bdf, 1'h1)
`STIMULI(5'h0f, 5'h08, 5'h09, 32'hc963a492, 1'h1)
`STIMULI(5'h0e, 5'h02, 5'h0a, 32'h76186bec, 1'h0)
`STIMULI(5'h02, 5'h03, 5'h0b, 32'h923adc24, 1'h1)
`STIMULI(5'h17, 5'h1f, 5'h0c, 32'hdb751eb6, 1'h0)
`STIMULI(5'h19, 5'h19, 5'h0d, 32'h04465108, 1'h1)
`STIMULI(5'h1c, 5'h0f, 5'h0e, 32'ha32d7646, 1'h0)
`STIMULI(5'h07, 5'h02, 5'h0f, 32'h4c41fb98, 1'h1)
`STIMULI(5'h00, 5'h0a, 5'h10, 32'hfb505ef6, 1'h0)
`STIMULI(5'h03, 5'h07, 5'h11, 32'hbf76227e, 1'h1)
`STIMULI(5'h17, 5'h02, 5'h12, 32'h9bcbfe37, 1'h0)
`STIMULI(5'h0f, 5'h17, 5'h13, 32'h44dbfb89, 1'h1)
`STIMULI(5'h1a, 5'h1e, 5'h14, 32'h3dc6dd7b, 1'h0)
`STIMULI(5'h19, 5'h13, 5'h15, 32'hd3a53ea7, 1'h1)
`STIMULI(5'h03, 5'h1e, 5'h16, 32'h1757fb2e, 1'h0)
`STIMULI(5'h1e, 5'h07, 5'h17, 32'h01cedd03, 1'h1)
`STIMULI(5'h16, 5'h0c, 5'h18, 32'h6165f1c2, 1'h0)
`STIMULI(5'h1d, 5'h05, 5'h19, 32'h4a268b94, 1'h0)
`STIMULI(5'h16, 5'h03, 5'h1a, 32'he9351ad2, 1'h0)
`STIMULI(5'h07, 5'h12, 5'h1b, 32'h67eb6bcf, 1'h1)
`STIMULI(5'h11, 5'h06, 5'h1c, 32'hfcecacf9, 1'h0)
`STIMULI(5'h18, 5'h0c, 5'h1d, 32'h16f1a92d, 1'h0)
`STIMULI(5'h00, 5'h0a, 5'h1e, 32'h921ad424, 1'h1)
`STIMULI(5'h1b, 5'h18, 5'h1f, 32'h61f123c3, 1'h1)
`STIMULI(5'h15, 5'h1e, 5'h00, 32'hc6ffe28d, 1'h1)
`STIMULI(5'h05, 5'h1b, 5'h01, 32'h9d66fe3a, 1'h1)
`STIMULI(5'h00, 5'h14, 5'h02, 32'hc3285e86, 1'h1)
`STIMULI(5'h1a, 5'h00, 5'h03, 32'hec324cd8, 1'h0)
`STIMULI(5'h17, 5'h0a, 5'h04, 32'hf19e2ae3, 1'h1)
`STIMULI(5'h18, 5'h13, 5'h05, 32'he3d3aec7, 1'h1)
`STIMULI(5'h11, 5'h0a, 5'h06, 32'h86b8a80d, 1'h0)
`STIMULI(5'h1e, 5'h16, 5'h07, 32'h48f7eb91, 1'h1)
`STIMULI(5'h01, 5'h13, 5'h08, 32'had53d45a, 1'h0)
`STIMULI(5'h13, 5'h18, 5'h09, 32'h19b59d33, 1'h1)
`STIMULI(5'h11, 5'h05, 5'h0a, 32'h82f66805, 1'h1)
`STIMULI(5'h1b, 5'h15, 5'h0b, 32'he1a5c2c3, 1'h1)
`STIMULI(5'h09, 5'h15, 5'h0c, 32'ha82ef650, 1'h1)
`STIMULI(5'h03, 5'h0d, 5'h0d, 32'hd4bf6ca9, 1'h1)
`STIMULI(5'h11, 5'h13, 5'h0e, 32'h8a301014, 1'h0)
`STIMULI(5'h0c, 5'h12, 5'h0f, 32'h189e5731, 1'h1)
`STIMULI(5'h0e, 5'h00, 5'h10, 32'h1c736538, 1'h0)
`STIMULI(5'h17, 5'h1e, 5'h11, 32'h289c8551, 1'h1)
`STIMULI(5'h13, 5'h19, 5'h12, 32'h6cebd9d9, 1'h1)
`STIMULI(5'h1f, 5'h0d, 5'h13, 32'h0fe6ed1f, 1'h1)
`STIMULI(5'h04, 5'h15, 5'h14, 32'hc30eb286, 1'h1)
`STIMULI(5'h1d, 5'h0b, 5'h15, 32'h7d7509fa, 1'h0)
`STIMULI(5'h16, 5'h1d, 5'h16, 32'hc1bbb283, 1'h1)
`STIMULI(5'h02, 5'h10, 5'h17, 32'h288b8551, 1'h1)
`STIMULI(5'h1a, 5'h19, 5'h18, 32'hbdcc347b, 1'h1)
`STIMULI(5'h1a, 5'h09, 5'h19, 32'hc931da92, 1'h1)
`STIMULI(5'h0b, 5'h1e, 5'h1a, 32'h16d1512d, 1'h0)
`STIMULI(5'h1b, 5'h02, 5'h1b, 32'hbec2e87d, 1'h0)
`STIMULI(5'h06, 5'h0c, 5'h1c, 32'h4d48fd9a, 1'h0)
`STIMULI(5'h1c, 5'h1a, 5'h1d, 32'h8f809e1f, 1'h1)
`STIMULI(5'h04, 5'h09, 5'h1e, 32'hc1522882, 1'h1)
`STIMULI(5'h1b, 5'h15, 5'h1f, 32'h66d297cd, 1'h0)
`STIMULI(5'h16, 5'h0f, 5'h00, 32'he6a7e2cd, 1'h0)
`STIMULI(5'h02, 5'h0b, 5'h01, 32'hcc97b899, 1'h0)
`STIMULI(5'h1c, 5'h02, 5'h02, 32'h3e6b6f7c, 1'h1)
`STIMULI(5'h1e, 5'h02, 5'h03, 32'haeb2d65d, 1'h1)
`STIMULI(5'h12, 5'h1a, 5'h04, 32'hfd0576fa, 1'h1)
`STIMULI(5'h1c, 5'h13, 5'h05, 32'haeba4e5d, 1'h0)
`STIMULI(5'h0b, 5'h04, 5'h06, 32'hda2616b4, 1'h0)
`STIMULI(5'h00, 5'h0b, 5'h07, 32'h2872ab50, 1'h1)
`STIMULI(5'h1b, 5'h0d, 5'h08, 32'h92ac0e25, 1'h0)
`STIMULI(5'h1d, 5'h0f, 5'h09, 32'hc27c4284, 1'h0)
`STIMULI(5'h18, 5'h03, 5'h0a, 32'h0ffad51f, 1'h0)
`STIMULI(5'h0f, 5'h10, 5'h0b, 32'h415bd982, 1'h0)
`STIMULI(5'h0c, 5'h0b, 5'h0c, 32'h6607bfcc, 1'h0)
`STIMULI(5'h13, 5'h0c, 5'h0d, 32'hf5c63aeb, 1'h0)
`STIMULI(5'h1c, 5'h0f, 5'h0e, 32'hd9261cb2, 1'h1)
`STIMULI(5'h17, 5'h0d, 5'h0f, 32'h29d6e353, 1'h1)
`STIMULI(5'h1c, 5'h15, 5'h10, 32'h4e5a5b9c, 1'h0)
`STIMULI(5'h1f, 5'h1b, 5'h11, 32'h9599982b, 1'h0)
`STIMULI(5'h01, 5'h0b, 5'h12, 32'hdcbc22b9, 1'h0)
`STIMULI(5'h0b, 5'h14, 5'h13, 32'hd20f0ea4, 1'h0)
`STIMULI(5'h00, 5'h05, 5'h14, 32'h1c2f7738, 1'h0)
`STIMULI(5'h06, 5'h09, 5'h15, 32'h2a948155, 1'h1)
`STIMULI(5'h07, 5'h00, 5'h16, 32'h357cd96a, 1'h1)
`STIMULI(5'h0d, 5'h13, 5'h17, 32'hbf565c7e, 1'h1)
`STIMULI(5'h14, 5'h1a, 5'h18, 32'h11906723, 1'h1)
`STIMULI(5'h0c, 5'h0e, 5'h19, 32'hd835d8b0, 1'h1)
`STIMULI(5'h18, 5'h01, 5'h1a, 32'h4167f782, 1'h0)
`STIMULI(5'h03, 5'h19, 5'h1b, 32'h3e49977c, 1'h0)
`STIMULI(5'h1d, 5'h12, 5'h1c, 32'hc5f83c8b, 1'h0)
`STIMULI(5'h00, 5'h0d, 5'h1d, 32'ha2e14245, 1'h0)
`STIMULI(5'h0f, 5'h0a, 5'h1e, 32'haf10ec5e, 1'h1)
`STIMULI(5'h03, 5'h12, 5'h1f, 32'h35b43b6b, 1'h1)
`STIMULI(5'h19, 5'h02, 5'h00, 32'h0a07d114, 1'h1)
`STIMULI(5'h1b, 5'h04, 5'h01, 32'hc0a32481, 1'h1)
`STIMULI(5'h01, 5'h1e, 5'h02, 32'hbcb2f079, 1'h1)
`STIMULI(5'h15, 5'h07, 5'h03, 32'h9e34903c, 1'h0)
`STIMULI(5'h1a, 5'h10, 5'h04, 32'h1ef9b33d, 1'h0)
`STIMULI(5'h05, 5'h0e, 5'h05, 32'hd8b4a0b1, 1'h0)
`STIMULI(5'h05, 5'h04, 5'h06, 32'h5d04f7ba, 1'h1)
`STIMULI(5'h1d, 5'h10, 5'h07, 32'h629f9bc5, 1'h0)
`STIMULI(5'h0a, 5'h1e, 5'h08, 32'h55d639ab, 1'h0)
`STIMULI(5'h1b, 5'h15, 5'h09, 32'hd5bf9aab, 1'h0)
`STIMULI(5'h12, 5'h03, 5'h0a, 32'hb5cdb26b, 1'h1)
`STIMULI(5'h0d, 5'h19, 5'h0b, 32'h2d251f5a, 1'h0)
`STIMULI(5'h18, 5'h1e, 5'h0c, 32'hea6778d4, 1'h1)
`STIMULI(5'h09, 5'h00, 5'h0d, 32'haee2b85d, 1'h1)
`STIMULI(5'h04, 5'h06, 5'h0e, 32'h2c379958, 1'h1)
`STIMULI(5'h0d, 5'h04, 5'h0f, 32'h65339fca, 1'h1)
`STIMULI(5'h06, 5'h0d, 5'h10, 32'haded425b, 1'h0)
`STIMULI(5'h19, 5'h19, 5'h11, 32'h4b755d96, 1'h0)
`STIMULI(5'h15, 5'h0d, 5'h12, 32'hf2e4dce5, 1'h0)
`STIMULI(5'h1f, 5'h16, 5'h13, 32'h621c61c4, 1'h1)
`STIMULI(5'h1c, 5'h06, 5'h14, 32'hd5912aab, 1'h1)
`STIMULI(5'h02, 5'h0c, 5'h15, 32'h658babcb, 1'h1)
`STIMULI(5'h03, 5'h18, 5'h16, 32'hcdc3709b, 1'h0)
`STIMULI(5'h03, 5'h05, 5'h17, 32'h9677662c, 1'h0)
`STIMULI(5'h17, 5'h11, 5'h18, 32'h009a8901, 1'h0)
`STIMULI(5'h02, 5'h05, 5'h19, 32'h0f3a891e, 1'h0)
`STIMULI(5'h17, 5'h0d, 5'h1a, 32'h7fa10dff, 1'h0)
`STIMULI(5'h08, 5'h0b, 5'h1b, 32'h38477570, 1'h1)
`STIMULI(5'h19, 5'h0e, 5'h1c, 32'h4a626f94, 1'h1)
`STIMULI(5'h1f, 5'h1c, 5'h1d, 32'h3e9b997d, 1'h1)
`STIMULI(5'h14, 5'h0f, 5'h1e, 32'h157f212a, 1'h0)
`STIMULI(5'h16, 5'h0d, 5'h1f, 32'ha9de0e53, 1'h0)
`STIMULI(5'h06, 5'h15, 5'h00, 32'hfc07aef8, 1'h0)
`STIMULI(5'h0c, 5'h0d, 5'h01, 32'h84913e09, 1'h1)
`STIMULI(5'h0e, 5'h19, 5'h02, 32'h03a6e307, 1'h0)
`STIMULI(5'h07, 5'h07, 5'h03, 32'ha77f7a4e, 1'h1)
`STIMULI(5'h0c, 5'h02, 5'h04, 32'h31e2e163, 1'h0)
`STIMULI(5'h1e, 5'h0f, 5'h05, 32'hd24aa0a4, 1'h1)
`STIMULI(5'h1b, 5'h18, 5'h06, 32'hc87d4690, 1'h1)
`STIMULI(5'h13, 5'h0a, 5'h07, 32'hfdc6bcfb, 1'h1)
`STIMULI(5'h0c, 5'h02, 5'h08, 32'h88ba5411, 1'h1)
`STIMULI(5'h19, 5'h08, 5'h09, 32'hf187a0e3, 1'h0)
`STIMULI(5'h02, 5'h02, 5'h0a, 32'h89170012, 1'h1)
`STIMULI(5'h1a, 5'h0f, 5'h0b, 32'h4cc99599, 1'h1)
`STIMULI(5'h1c, 5'h01, 5'h0c, 32'ha6b6204d, 1'h0)
`STIMULI(5'h1e, 5'h0c, 5'h0d, 32'h139ce527, 1'h0)
`STIMULI(5'h09, 5'h17, 5'h0e, 32'hdb8c84b7, 1'h1)
`STIMULI(5'h0b, 5'h01, 5'h0f, 32'h1bfc8b37, 1'h0)
`STIMULI(5'h00, 5'h01, 5'h10, 32'h34141968, 1'h0)
`STIMULI(5'h1c, 5'h0e, 5'h11, 32'h9b37ce36, 1'h0)
`STIMULI(5'h18, 5'h0b, 5'h12, 32'hb30e0466, 1'h1)
`STIMULI(5'h1f, 5'h17, 5'h13, 32'h42d6e385, 1'h0)
`STIMULI(5'h1f, 5'h0c, 5'h14, 32'h979bd02f, 1'h0)
`STIMULI(5'h17, 5'h0c, 5'h15, 32'h04e28309, 1'h1)
`STIMULI(5'h0f, 5'h11, 5'h16, 32'h21b77943, 1'h0)
`STIMULI(5'h1f, 5'h16, 5'h17, 32'h6a369fd4, 1'h1)
`STIMULI(5'h0c, 5'h16, 5'h18, 32'h8ad29a15, 1'h1)
`STIMULI(5'h1f, 5'h19, 5'h19, 32'h9247e624, 1'h1)
`STIMULI(5'h18, 5'h1d, 5'h1a, 32'h642491c8, 1'h0)
`STIMULI(5'h0e, 5'h02, 5'h1b, 32'h2a848355, 1'h1)
`STIMULI(5'h18, 5'h12, 5'h1c, 32'h59ef8fb3, 1'h0)
`STIMULI(5'h0e, 5'h12, 5'h1d, 32'h1c379d38, 1'h1)
`STIMULI(5'h1f, 5'h10, 5'h1e, 32'h6ac4c5d5, 1'h1)
`STIMULI(5'h0c, 5'h1b, 5'h1f, 32'h0a981315, 1'h1)
`STIMULI(5'h1e, 5'h1f, 5'h00, 32'h638f7fc7, 1'h0)
`STIMULI(5'h06, 5'h08, 5'h01, 32'h2f6a0b5e, 1'h0)
`STIMULI(5'h19, 5'h1a, 5'h02, 32'hd4ef44a9, 1'h0)
`STIMULI(5'h14, 5'h12, 5'h03, 32'h635b95c6, 1'h0)
`STIMULI(5'h18, 5'h1d, 5'h04, 32'h2c28fd58, 1'h0)
`STIMULI(5'h08, 5'h1a, 5'h05, 32'h580453b0, 1'h0)
`STIMULI(5'h1f, 5'h07, 5'h06, 32'h11b70723, 1'h0)
`STIMULI(5'h1a, 5'h14, 5'h07, 32'hec300cd8, 1'h1)
`STIMULI(5'h15, 5'h0d, 5'h08, 32'h19405f32, 1'h1)
`STIMULI(5'h15, 5'h1e, 5'h09, 32'h3fdc597f, 1'h1)
`STIMULI(5'h07, 5'h16, 5'h0a, 32'h1a7ebf34, 1'h1)
`STIMULI(5'h16, 5'h07, 5'h0b, 32'h74113be8, 1'h1)
`STIMULI(5'h02, 5'h1e, 5'h0c, 32'ha85bb850, 1'h1)
`STIMULI(5'h01, 5'h07, 5'h0d, 32'h037cc306, 1'h1)
`STIMULI(5'h04, 5'h15, 5'h0e, 32'hfb4ce0f6, 1'h0)
`STIMULI(5'h07, 5'h03, 5'h0f, 32'h0b79a716, 1'h0)
`STIMULI(5'h14, 5'h04, 5'h10, 32'hb5b6de6b, 1'h1)
`STIMULI(5'h18, 5'h05, 5'h11, 32'he1e8f2c3, 1'h1)
`STIMULI(5'h0f, 5'h08, 5'h12, 32'h1cdf9f39, 1'h1)
`STIMULI(5'h08, 5'h15, 5'h13, 32'ha3069446, 1'h0)
`STIMULI(5'h07, 5'h1d, 5'h14, 32'h26b7654d, 1'h1)
`STIMULI(5'h04, 5'h18, 5'h15, 32'h2b210d56, 1'h1)
`STIMULI(5'h0b, 5'h0e, 5'h16, 32'h0480f109, 1'h0)
`STIMULI(5'h15, 5'h0d, 5'h17, 32'he2dc06c5, 1'h1)
`STIMULI(5'h15, 5'h1a, 5'h18, 32'h0c209f18, 1'h0)
`STIMULI(5'h01, 5'h0c, 5'h19, 32'h1165f722, 1'h1)
`STIMULI(5'h05, 5'h01, 5'h1a, 32'hfd9a86fb, 1'h1)
`STIMULI(5'h0e, 5'h1f, 5'h1b, 32'hbec8c07d, 1'h1)
`STIMULI(5'h0d, 5'h03, 5'h1c, 32'h10079f20, 1'h0)
`STIMULI(5'h18, 5'h17, 5'h1d, 32'hc13d5282, 1'h1)
`STIMULI(5'h15, 5'h1f, 5'h1e, 32'he109d8c2, 1'h0)
`STIMULI(5'h18, 5'h08, 5'h1f, 32'h0b2a4716, 1'h1)
`STIMULI(5'h17, 5'h0e, 5'h00, 32'hc3873c87, 1'h1)
`STIMULI(5'h14, 5'h0c, 5'h01, 32'he43584c8, 1'h0)
`STIMULI(5'h12, 5'h01, 5'h02, 32'hee3416dc, 1'h0)
`STIMULI(5'h15, 5'h0f, 5'h03, 32'h1690df2d, 1'h0)
`STIMULI(5'h0a, 5'h06, 5'h04, 32'h20340940, 1'h1)
`STIMULI(5'h1c, 5'h0a, 5'h05, 32'h7269b3e4, 1'h0)
`STIMULI(5'h19, 5'h10, 5'h06, 32'h69da37d3, 1'h0)
`STIMULI(5'h01, 5'h00, 5'h07, 32'h0c238d18, 1'h0)
`STIMULI(5'h13, 5'h0b, 5'h08, 32'h515059a2, 1'h0)
`STIMULI(5'h0a, 5'h06, 5'h09, 32'h76c5c1ed, 1'h0)
`STIMULI(5'h15, 5'h0d, 5'h0a, 32'h76aceded, 1'h1)
`STIMULI(5'h17, 5'h0f, 5'h0b, 32'ha2c41045, 1'h0)
`STIMULI(5'h0a, 5'h1a, 5'h0c, 32'h98c04231, 1'h0)
`STIMULI(5'h1b, 5'h05, 5'h0d, 32'h2a0a4f54, 1'h0)
`STIMULI(5'h04, 5'h0d, 5'h0e, 32'h5ba0abb7, 1'h1)
`STIMULI(5'h0d, 5'h04, 5'h0f, 32'h5cf2f3b9, 1'h0)
`STIMULI(5'h06, 5'h01, 5'h10, 32'he3bd96c7, 1'h1)
`STIMULI(5'h12, 5'h03, 5'h11, 32'h8890c411, 1'h1)
`STIMULI(5'h13, 5'h00, 5'h12, 32'h2c01a958, 1'h0)
`STIMULI(5'h0e, 5'h02, 5'h13, 32'h5d7377ba, 1'h1)
`STIMULI(5'h0c, 5'h1d, 5'h14, 32'h634be9c6, 1'h0)
`STIMULI(5'h1d, 5'h19, 5'h15, 32'h46cf478d, 1'h0)
`STIMULI(5'h0d, 5'h09, 5'h16, 32'h8547d80a, 1'h0)
`STIMULI(5'h0f, 5'h09, 5'h17, 32'h94af9e29, 1'h0)
`STIMULI(5'h0a, 5'h04, 5'h18, 32'h3c6c9178, 1'h1)
`STIMULI(5'h1c, 5'h1a, 5'h19, 32'hc89cb491, 1'h1)
`STIMULI(5'h1f, 5'h04, 5'h1a, 32'hd6aaecad, 1'h1)
`STIMULI(5'h1a, 5'h1d, 5'h1b, 32'hcadc2e95, 1'h1)
`STIMULI(5'h06, 5'h01, 5'h1c, 32'h2412a148, 1'h0)
`STIMULI(5'h00, 5'h08, 5'h1d, 32'h7f34b9fe, 1'h0)
`STIMULI(5'h11, 5'h03, 5'h1e, 32'h66765bcc, 1'h1)
`STIMULI(5'h02, 5'h19, 5'h1f, 32'hcadcaa95, 1'h0)
`STIMULI(5'h02, 5'h09, 5'h00, 32'h7ad6ebf5, 1'h1)
`STIMULI(5'h1a, 5'h0c, 5'h01, 32'hd1fbb0a3, 1'h1)
`STIMULI(5'h1f, 5'h07, 5'h02, 32'h091d5712, 1'h1)
`STIMULI(5'h1b, 5'h00, 5'h03, 32'hb1e75863, 1'h0)
`STIMULI(5'h05, 5'h1b, 5'h04, 32'h3c6c0778, 1'h1)
`STIMULI(5'h0d, 5'h13, 5'h05, 32'h7602c5ec, 1'h1)
`STIMULI(5'h0d, 5'h0a, 5'h06, 32'h3e0ed77c, 1'h0)
`STIMULI(5'h10, 5'h1a, 5'h07, 32'h27e93d4f, 1'h1)
`STIMULI(5'h0c, 5'h01, 5'h08, 32'hd6d244ad, 1'h1)
`STIMULI(5'h07, 5'h06, 5'h09, 32'hd84bd6b0, 1'h1)
`STIMULI(5'h19, 5'h0c, 5'h0a, 32'h2649894c, 1'h1)
`STIMULI(5'h0a, 5'h0f, 5'h0b, 32'h04aa1709, 1'h0)
`STIMULI(5'h0d, 5'h10, 5'h0c, 32'hbd4bba7a, 1'h0)
`STIMULI(5'h0a, 5'h0d, 5'h0d, 32'hfecd8cfd, 1'h0)
`STIMULI(5'h11, 5'h05, 5'h0e, 32'h88afe611, 1'h1)
`STIMULI(5'h03, 5'h15, 5'h0f, 32'ha5b06e4b, 1'h1)
`STIMULI(5'h13, 5'h19, 5'h10, 32'h4b103d96, 1'h1)
`STIMULI(5'h0a, 5'h05, 5'h11, 32'h04374908, 1'h0)
`STIMULI(5'h19, 5'h06, 5'h12, 32'hd81c22b0, 1'h1)
`STIMULI(5'h1d, 5'h0b, 5'h13, 32'hf8e588f1, 1'h0)
`STIMULI(5'h1b, 5'h04, 5'h14, 32'h49c15f93, 1'h0)
`STIMULI(5'h10, 5'h0d, 5'h15, 32'h12752f24, 1'h1)
`STIMULI(5'h01, 5'h16, 5'h16, 32'hef342ede, 1'h1)
`STIMULI(5'h12, 5'h01, 5'h17, 32'hfff966ff, 1'h0)
`STIMULI(5'h1e, 5'h15, 5'h18, 32'h2f9e735f, 1'h0)
`STIMULI(5'h1e, 5'h14, 5'h19, 32'h7ff425ff, 1'h1)
`STIMULI(5'h1f, 5'h07, 5'h1a, 32'hf5fdc2eb, 1'h0)
`STIMULI(5'h1e, 5'h0d, 5'h1b, 32'h5086cda1, 1'h1)
`STIMULI(5'h07, 5'h03, 5'h1c, 32'he97890d2, 1'h0)
`STIMULI(5'h04, 5'h19, 5'h1d, 32'h73a5cde7, 1'h1)
`STIMULI(5'h08, 5'h1e, 5'h1e, 32'ha5324e4a, 1'h1)
`STIMULI(5'h0c, 5'h0c, 5'h1f, 32'hd4f740a9, 1'h0)
`STIMULI(5'h05, 5'h0d, 5'h00, 32'hc4668888, 1'h1)
`STIMULI(5'h13, 5'h0e, 5'h01, 32'h33c48d67, 1'h1)
`STIMULI(5'h00, 5'h1a, 5'h02, 32'hdb5308b6, 1'h1)
`STIMULI(5'h0c, 5'h1b, 5'h03, 32'hd22702a4, 1'h0)
`STIMULI(5'h02, 5'h10, 5'h04, 32'hcb38f296, 1'h0)
`STIMULI(5'h05, 5'h00, 5'h05, 32'h03578506, 1'h0)
`STIMULI(5'h14, 5'h04, 5'h06, 32'h377ce56e, 1'h1)
`STIMULI(5'h05, 5'h04, 5'h07, 32'hf5c91ceb, 1'h0)
`STIMULI(5'h1e, 5'h0b, 5'h08, 32'habae1e57, 1'h0)
`STIMULI(5'h16, 5'h1d, 5'h09, 32'h32769f64, 1'h1)
`STIMULI(5'h18, 5'h12, 5'h0a, 32'h2dfc975b, 1'h0)
`STIMULI(5'h16, 5'h03, 5'h0b, 32'hf18b4ce3, 1'h0)
`STIMULI(5'h1b, 5'h13, 5'h0c, 32'hf76622ee, 1'h1)
`STIMULI(5'h07, 5'h03, 5'h0d, 32'hc54e788a, 1'h0)
`STIMULI(5'h0d, 5'h19, 5'h0e, 32'hcaa29295, 1'h0)
`STIMULI(5'h07, 5'h1f, 5'h0f, 32'he6fa1ccd, 1'h1)
`STIMULI(5'h0d, 5'h07, 5'h10, 32'h5496d3a9, 1'h1)
`STIMULI(5'h17, 5'h00, 5'h11, 32'hd5e47aab, 1'h0)
`STIMULI(5'h0c, 5'h07, 5'h12, 32'h14d70d29, 1'h0)
`STIMULI(5'h19, 5'h15, 5'h13, 32'ha824ca50, 1'h0)
`STIMULI(5'h1c, 5'h04, 5'h14, 32'hf27fc2e4, 1'h1)
`STIMULI(5'h04, 5'h0c, 5'h15, 32'h949ac829, 1'h1)
`STIMULI(5'h0f, 5'h1e, 5'h16, 32'hc96df692, 1'h0)
`STIMULI(5'h18, 5'h04, 5'h17, 32'h91015e22, 1'h1)
`STIMULI(5'h1b, 5'h05, 5'h18, 32'h559e47ab, 1'h1)
`STIMULI(5'h0a, 5'h06, 5'h19, 32'h8b744216, 1'h0)
`STIMULI(5'h15, 5'h05, 5'h1a, 32'hde3b08bc, 1'h1)
`STIMULI(5'h1b, 5'h1a, 5'h1b, 32'h7d909bfb, 1'h0)
`STIMULI(5'h0d, 5'h19, 5'h1c, 32'h4fa1719f, 1'h1)
`STIMULI(5'h16, 5'h1a, 5'h1d, 32'h88189210, 1'h1)
`STIMULI(5'h06, 5'h08, 5'h1e, 32'h0365b306, 1'h1)
`STIMULI(5'h0f, 5'h16, 5'h1f, 32'h20c20541, 1'h0)
`STIMULI(5'h01, 5'h11, 5'h00, 32'hb71e186e, 1'h1)
`STIMULI(5'h10, 5'h14, 5'h01, 32'h509817a1, 1'h1)
`STIMULI(5'h0d, 5'h02, 5'h02, 32'h167d2b2c, 1'h0)
`STIMULI(5'h0a, 5'h11, 5'h03, 32'hc017de80, 1'h1)
`STIMULI(5'h15, 5'h14, 5'h04, 32'h3302cf66, 1'h0)
`STIMULI(5'h05, 5'h15, 5'h05, 32'h06eff70d, 1'h1)
`STIMULI(5'h00, 5'h04, 5'h06, 32'h3b4c6576, 1'h0)
`STIMULI(5'h19, 5'h1a, 5'h07, 32'h180b2d30, 1'h0)
`STIMULI(5'h1d, 5'h1d, 5'h08, 32'h2dcbe95b, 1'h1)
`STIMULI(5'h18, 5'h02, 5'h09, 32'hdf4e14be, 1'h1)
`STIMULI(5'h10, 5'h14, 5'h0a, 32'h0e6e151c, 1'h1)
`STIMULI(5'h1a, 5'h01, 5'h0b, 32'hed2fb4da, 1'h1)
`STIMULI(5'h1d, 5'h0e, 5'h0c, 32'hc4777a88, 1'h0)
`STIMULI(5'h01, 5'h00, 5'h0d, 32'h8d15161a, 1'h0)
`STIMULI(5'h0e, 5'h1e, 5'h0e, 32'h25a0af4b, 1'h1)
`STIMULI(5'h0d, 5'h03, 5'h0f, 32'h8e17f81c, 1'h1)
`STIMULI(5'h00, 5'h1d, 5'h10, 32'h4539598a, 1'h1)
`STIMULI(5'h07, 5'h00, 5'h11, 32'h8aa05e15, 1'h0)
`STIMULI(5'h0d, 5'h07, 5'h12, 32'hd1da66a3, 1'h0)
`STIMULI(5'h1f, 5'h1a, 5'h13, 32'h49f93d93, 1'h1)
`STIMULI(5'h0c, 5'h06, 5'h14, 32'h91ef1623, 1'h1)
`STIMULI(5'h17, 5'h06, 5'h15, 32'h1fc8113f, 1'h0)
`STIMULI(5'h15, 5'h06, 5'h16, 32'hd71d2eae, 1'h1)
`STIMULI(5'h15, 5'h1a, 5'h17, 32'ha00f8640, 1'h1)
`STIMULI(5'h01, 5'h04, 5'h18, 32'h7a5409f4, 1'h1)
`STIMULI(5'h1f, 5'h12, 5'h19, 32'hcb251296, 1'h1)
`STIMULI(5'h0c, 5'h0f, 5'h1a, 32'h8e0abc1c, 1'h0)
`STIMULI(5'h0b, 5'h06, 5'h1b, 32'habc19857, 1'h1)
`STIMULI(5'h0b, 5'h0b, 5'h1c, 32'he1f542c3, 1'h0)
`STIMULI(5'h02, 5'h0f, 5'h1d, 32'h721507e4, 1'h0)
`STIMULI(5'h0e, 5'h12, 5'h1e, 32'ha3388646, 1'h0)
`STIMULI(5'h1c, 5'h03, 5'h1f, 32'h1184f923, 1'h1)
`STIMULI(5'h0d, 5'h04, 5'h00, 32'h45e5978b, 1'h0)
`STIMULI(5'h1d, 5'h16, 5'h01, 32'h7b7e53f6, 1'h0)
`STIMULI(5'h13, 5'h00, 5'h02, 32'h6843bdd0, 1'h1)
`STIMULI(5'h0d, 5'h0a, 5'h03, 32'h7081e9e1, 1'h0)
`STIMULI(5'h08, 5'h0c, 5'h04, 32'hf6319aec, 1'h1)
`STIMULI(5'h07, 5'h0e, 5'h05, 32'hb9541872, 1'h0)
`STIMULI(5'h1d, 5'h09, 5'h06, 32'h6aa555d5, 1'h0)
`STIMULI(5'h1a, 5'h0f, 5'h07, 32'h1cf76d39, 1'h0)
`STIMULI(5'h18, 5'h04, 5'h08, 32'h1713a52e, 1'h1)
`STIMULI(5'h04, 5'h03, 5'h09, 32'hc4da3c89, 1'h0)
`STIMULI(5'h15, 5'h01, 5'h0a, 32'hc4460288, 1'h0)
`STIMULI(5'h0c, 5'h19, 5'h0b, 32'ha75f4a4e, 1'h0)
`STIMULI(5'h14, 5'h05, 5'h0c, 32'h3de7c57b, 1'h1)
`STIMULI(5'h01, 5'h14, 5'h0d, 32'h31a96363, 1'h1)
`STIMULI(5'h05, 5'h00, 5'h0e, 32'h59d23bb3, 1'h0)
`STIMULI(5'h04, 5'h1b, 5'h0f, 32'h745205e8, 1'h1)
`STIMULI(5'h10, 5'h06, 5'h10, 32'h3ddfd17b, 1'h1)
`STIMULI(5'h02, 5'h09, 5'h11, 32'hbb72f076, 1'h0)
`STIMULI(5'h1a, 5'h01, 5'h12, 32'hface2ef5, 1'h0)
`STIMULI(5'h03, 5'h0f, 5'h13, 32'h692adfd2, 1'h0)
`STIMULI(5'h02, 5'h0b, 5'h14, 32'h78775df0, 1'h1)
`STIMULI(5'h1d, 5'h02, 5'h15, 32'h52850ba5, 1'h0)
`STIMULI(5'h08, 5'h07, 5'h16, 32'h1769d72e, 1'h1)
`STIMULI(5'h14, 5'h00, 5'h17, 32'h716bdfe2, 1'h1)
`STIMULI(5'h0a, 5'h1c, 5'h18, 32'hc5a7ba8b, 1'h0)
`STIMULI(5'h10, 5'h12, 5'h19, 32'hab0e9256, 1'h1)
`STIMULI(5'h03, 5'h0f, 5'h1a, 32'h8014e200, 1'h0)
`STIMULI(5'h02, 5'h0b, 5'h1b, 32'h60e1c7c1, 1'h1)
`STIMULI(5'h10, 5'h16, 5'h1c, 32'hc7dc028f, 1'h0)
`STIMULI(5'h0d, 5'h15, 5'h1d, 32'hb3232c66, 1'h1)
`STIMULI(5'h1e, 5'h06, 5'h1e, 32'h62d2cbc5, 1'h0)
`STIMULI(5'h1d, 5'h1a, 5'h1f, 32'h76881ded, 1'h1)
`STIMULI(5'h18, 5'h0b, 5'h00, 32'h3fa5057f, 1'h1)
`STIMULI(5'h1c, 5'h05, 5'h01, 32'h137f3d26, 1'h0)
`STIMULI(5'h1a, 5'h0b, 5'h02, 32'h7a4ebff4, 1'h1)
`STIMULI(5'h06, 5'h07, 5'h03, 32'h842d2208, 1'h1)
`STIMULI(5'h1e, 5'h15, 5'h04, 32'hb32d5866, 1'h0)
`STIMULI(5'h1d, 5'h1d, 5'h05, 32'h9f0be83e, 1'h1)
`STIMULI(5'h0a, 5'h0b, 5'h06, 32'h22afb545, 1'h0)
`STIMULI(5'h10, 5'h0e, 5'h07, 32'h7ed5ddfd, 1'h1)
`STIMULI(5'h14, 5'h04, 5'h08, 32'h7d6d4ffa, 1'h0)
`STIMULI(5'h0d, 5'h07, 5'h09, 32'h552313aa, 1'h0)
`STIMULI(5'h15, 5'h1d, 5'h0a, 32'hc82c6090, 1'h1)
`STIMULI(5'h1a, 5'h10, 5'h0b, 32'hfbe210f7, 1'h0)
`STIMULI(5'h17, 5'h13, 5'h0c, 32'h191efd32, 1'h0)
`STIMULI(5'h05, 5'h0b, 5'h0d, 32'h5a9361b5, 1'h0)
`STIMULI(5'h19, 5'h06, 5'h0e, 32'he35f34c6, 1'h1)
`STIMULI(5'h10, 5'h17, 5'h0f, 32'hdef040bd, 1'h0)
`STIMULI(5'h18, 5'h03, 5'h10, 32'h3b723776, 1'h0)
`STIMULI(5'h05, 5'h18, 5'h11, 32'h0d64351a, 1'h0)
`STIMULI(5'h03, 5'h09, 5'h12, 32'h775a69ee, 1'h0)
`STIMULI(5'h12, 5'h01, 5'h13, 32'h3c81b179, 1'h0)
`STIMULI(5'h0e, 5'h0c, 5'h14, 32'h12809125, 1'h0)
`STIMULI(5'h05, 5'h00, 5'h15, 32'h1759b32e, 1'h0)
`STIMULI(5'h17, 5'h14, 5'h16, 32'hc57bee8a, 1'h1)
`STIMULI(5'h19, 5'h10, 5'h17, 32'h355e676a, 1'h1)
`STIMULI(5'h09, 5'h0c, 5'h18, 32'hbb815e77, 1'h1)
`STIMULI(5'h0b, 5'h19, 5'h19, 32'h2338c146, 1'h0)
`STIMULI(5'h14, 5'h07, 5'h1a, 32'hab017856, 1'h0)
`STIMULI(5'h08, 5'h1b, 5'h1b, 32'h4eb9259d, 1'h1)
`STIMULI(5'h1e, 5'h13, 5'h1c, 32'hc4bdb289, 1'h0)
`STIMULI(5'h12, 5'h04, 5'h1d, 32'h98cb0031, 1'h1)
`STIMULI(5'h08, 5'h04, 5'h1e, 32'hdc5c7cb8, 1'h1)
`STIMULI(5'h13, 5'h16, 5'h1f, 32'h8b137016, 1'h1)
`STIMULI(5'h0a, 5'h05, 5'h00, 32'h4f44659e, 1'h1)
`STIMULI(5'h09, 5'h0a, 5'h01, 32'h83a2d807, 1'h1)
`STIMULI(5'h01, 5'h13, 5'h02, 32'hf24630e4, 1'h0)
`STIMULI(5'h1c, 5'h1e, 5'h03, 32'h47e18d8f, 1'h0)
`STIMULI(5'h11, 5'h03, 5'h04, 32'h245e0548, 1'h0)
`STIMULI(5'h10, 5'h10, 5'h05, 32'h889f6a11, 1'h0)
`STIMULI(5'h03, 5'h17, 5'h06, 32'hfc9384f9, 1'h0)
`STIMULI(5'h1a, 5'h19, 5'h07, 32'ha3ee7c47, 1'h1)
`STIMULI(5'h0f, 5'h19, 5'h08, 32'hd2c0e8a5, 1'h1)
`STIMULI(5'h1b, 5'h0c, 5'h09, 32'h8e309a1c, 1'h1)
`STIMULI(5'h14, 5'h06, 5'h0a, 32'h0ec92d1d, 1'h1)
`STIMULI(5'h0a, 5'h03, 5'h0b, 32'hf28006e5, 1'h0)
`STIMULI(5'h18, 5'h0b, 5'h0c, 32'ha785244f, 1'h0)
`STIMULI(5'h07, 5'h04, 5'h0d, 32'h7b5b0ff6, 1'h0)
`STIMULI(5'h0c, 5'h0a, 5'h0e, 32'hfa6fa0f4, 1'h1)
`STIMULI(5'h0e, 5'h01, 5'h0f, 32'h7f3aadfe, 1'h1)
`STIMULI(5'h0c, 5'h10, 5'h10, 32'h16d88d2d, 1'h1)
`STIMULI(5'h09, 5'h02, 5'h11, 32'h317c2962, 1'h0)
`STIMULI(5'h16, 5'h0b, 5'h12, 32'h2b271356, 1'h1)
`STIMULI(5'h0f, 5'h12, 5'h13, 32'ha6c5b24d, 1'h0)
`STIMULI(5'h14, 5'h1c, 5'h14, 32'he872b4d0, 1'h1)
`STIMULI(5'h15, 5'h18, 5'h15, 32'ha4ce0c49, 1'h0)
`STIMULI(5'h07, 5'h19, 5'h16, 32'h587b75b0, 1'h0)
`STIMULI(5'h1e, 5'h16, 5'h17, 32'h082f1f10, 1'h0)
`STIMULI(5'h05, 5'h0c, 5'h18, 32'h3bc8f177, 1'h0)
`STIMULI(5'h13, 5'h11, 5'h19, 32'hb7aba06f, 1'h0)
`STIMULI(5'h11, 5'h10, 5'h1a, 32'h81787e02, 1'h0)
`STIMULI(5'h02, 5'h00, 5'h1b, 32'h530fb3a6, 1'h0)
`STIMULI(5'h14, 5'h11, 5'h1c, 32'h38025570, 1'h0)
`STIMULI(5'h04, 5'h07, 5'h1d, 32'h3c948779, 1'h0)
`STIMULI(5'h19, 5'h04, 5'h1e, 32'h65fda1cb, 1'h0)
`STIMULI(5'h17, 5'h0d, 5'h1f, 32'hf66ef4ec, 1'h1)
`STIMULI(5'h03, 5'h09, 5'h00, 32'hfbabb2f7, 1'h1)
`STIMULI(5'h17, 5'h04, 5'h01, 32'h42f12385, 1'h1)
`STIMULI(5'h1f, 5'h00, 5'h02, 32'h71d211e3, 1'h1)
`STIMULI(5'h10, 5'h01, 5'h03, 32'hb4672668, 1'h1)
`STIMULI(5'h13, 5'h06, 5'h04, 32'h202ba140, 1'h0)
`STIMULI(5'h03, 5'h08, 5'h05, 32'h92969a25, 1'h0)
`STIMULI(5'h1a, 5'h15, 5'h06, 32'hcd78c29a, 1'h1)
`STIMULI(5'h0f, 5'h0d, 5'h07, 32'hde894cbd, 1'h1)
`STIMULI(5'h1e, 5'h18, 5'h08, 32'he4f674c9, 1'h0)
`STIMULI(5'h0e, 5'h08, 5'h09, 32'hfa0ad2f4, 1'h1)
`STIMULI(5'h10, 5'h14, 5'h0a, 32'h08c46b11, 1'h0)
`STIMULI(5'h1b, 5'h0a, 5'h0b, 32'hbf012c7e, 1'h1)
`STIMULI(5'h1f, 5'h19, 5'h0c, 32'hd6823ead, 1'h0)
`STIMULI(5'h15, 5'h1b, 5'h0d, 32'hd3886aa7, 1'h0)
`STIMULI(5'h14, 5'h03, 5'h0e, 32'h932b7c26, 1'h0)
`STIMULI(5'h14, 5'h19, 5'h0f, 32'h727949e4, 1'h0)
`STIMULI(5'h17, 5'h1e, 5'h10, 32'h84fad409, 1'h1)
`STIMULI(5'h1b, 5'h13, 5'h11, 32'he4c2cac9, 1'h1)
`STIMULI(5'h13, 5'h0b, 5'h12, 32'hf5dc2ceb, 1'h1)
`STIMULI(5'h18, 5'h00, 5'h13, 32'h36bee56d, 1'h0)
`STIMULI(5'h15, 5'h02, 5'h14, 32'h9eb5ca3d, 1'h1)
`STIMULI(5'h0a, 5'h18, 5'h15, 32'h7d6a17fa, 1'h1)
`STIMULI(5'h17, 5'h18, 5'h16, 32'h83906c07, 1'h0)
`STIMULI(5'h17, 5'h1b, 5'h17, 32'hf22606e4, 1'h1)
`STIMULI(5'h02, 5'h0d, 5'h18, 32'h82667204, 1'h0)
`STIMULI(5'h07, 5'h1e, 5'h19, 32'h786f2ff0, 1'h0)
`STIMULI(5'h01, 5'h1d, 5'h1a, 32'hf221f4e4, 1'h0)
`STIMULI(5'h08, 5'h1b, 5'h1b, 32'h77ad71ef, 1'h1)
`STIMULI(5'h05, 5'h18, 5'h1c, 32'h1d11e53a, 1'h1)
`STIMULI(5'h11, 5'h05, 5'h1d, 32'h8407ba08, 1'h0)
`STIMULI(5'h15, 5'h18, 5'h1e, 32'h11de3523, 1'h0)
`STIMULI(5'h1b, 5'h0c, 5'h1f, 32'hcbe2a897, 1'h1)
`STIMULI(5'h19, 5'h04, 5'h00, 32'ha7c2f04f, 1'h1)
`STIMULI(5'h0f, 5'h0d, 5'h01, 32'hd4721ea8, 1'h1)
`STIMULI(5'h03, 5'h11, 5'h02, 32'h969a622d, 1'h1)
`STIMULI(5'h1a, 5'h17, 5'h03, 32'h6e85f1dd, 1'h1)
`STIMULI(5'h10, 5'h01, 5'h04, 32'h98fe2e31, 1'h0)
`STIMULI(5'h10, 5'h02, 5'h05, 32'h25797d4a, 1'h0)
`STIMULI(5'h19, 5'h04, 5'h06, 32'ha687724d, 1'h0)
`STIMULI(5'h1f, 5'h1b, 5'h07, 32'h6cee4dd9, 1'h1)
`STIMULI(5'h0f, 5'h0d, 5'h08, 32'hddf5eebb, 1'h1)
`STIMULI(5'h00, 5'h0b, 5'h09, 32'haeb9b85d, 1'h0)
`STIMULI(5'h1e, 5'h12, 5'h0a, 32'ha2c61845, 1'h1)
`STIMULI(5'h03, 5'h11, 5'h0b, 32'hc12d8282, 1'h0)
`STIMULI(5'h0d, 5'h00, 5'h0c, 32'h2f7e475e, 1'h1)
`STIMULI(5'h18, 5'h1f, 5'h0d, 32'h6ea379dd, 1'h1)
`STIMULI(5'h02, 5'h1c, 5'h0e, 32'h5dbac9bb, 1'h1)
`STIMULI(5'h10, 5'h18, 5'h0f, 32'h41f41583, 1'h0)
`STIMULI(5'h1e, 5'h18, 5'h10, 32'h16c10b2d, 1'h1)
`STIMULI(5'h02, 5'h0f, 5'h11, 32'hf0401ee0, 1'h0)
`STIMULI(5'h18, 5'h04, 5'h12, 32'hb321b666, 1'h0)
`STIMULI(5'h1f, 5'h1f, 5'h13, 32'h2735474e, 1'h0)
`STIMULI(5'h06, 5'h01, 5'h14, 32'hf5b1ceeb, 1'h0)
`STIMULI(5'h1a, 5'h09, 5'h15, 32'h6fb5cfdf, 1'h1)
`STIMULI(5'h1d, 5'h0c, 5'h16, 32'h35e2d56b, 1'h0)
`STIMULI(5'h10, 5'h1e, 5'h17, 32'he78b1ecf, 1'h1)
`STIMULI(5'h19, 5'h17, 5'h18, 32'h2741e74e, 1'h1)
`STIMULI(5'h1b, 5'h19, 5'h19, 32'h018b6f03, 1'h0)
`STIMULI(5'h07, 5'h17, 5'h1a, 32'h67a5dbcf, 1'h0)
`STIMULI(5'h0d, 5'h08, 5'h1b, 32'hf25a5ee4, 1'h0)
`STIMULI(5'h1d, 5'h05, 5'h1c, 32'h0b546516, 1'h1)
`STIMULI(5'h1a, 5'h1b, 5'h1d, 32'h20aca141, 1'h1)
`STIMULI(5'h18, 5'h09, 5'h1e, 32'hae26385c, 1'h0)
`STIMULI(5'h08, 5'h18, 5'h1f, 32'h8ab68c15, 1'h1)
`STIMULI(5'h1e, 5'h1d, 5'h00, 32'h92722024, 1'h0)
`STIMULI(5'h15, 5'h15, 5'h01, 32'hc72dca8e, 1'h1)
`STIMULI(5'h15, 5'h1f, 5'h02, 32'hfa4724f4, 1'h1)
`STIMULI(5'h0a, 5'h01, 5'h03, 32'hc705ea8e, 1'h0)
`STIMULI(5'h09, 5'h12, 5'h04, 32'h9d3daa3a, 1'h1)
`STIMULI(5'h07, 5'h12, 5'h05, 32'hf5d00ceb, 1'h1)
`STIMULI(5'h01, 5'h1a, 5'h06, 32'hd4e792a9, 1'h1)
`STIMULI(5'h11, 5'h10, 5'h07, 32'h79657df2, 1'h0)
`STIMULI(5'h07, 5'h1c, 5'h08, 32'h43a75987, 1'h1)
`STIMULI(5'h01, 5'h1c, 5'h09, 32'h4e45519c, 1'h1)
`STIMULI(5'h0a, 5'h08, 5'h0a, 32'h4576378a, 1'h1)
`STIMULI(5'h10, 5'h00, 5'h0b, 32'h84cd0809, 1'h1)
`STIMULI(5'h1a, 5'h1b, 5'h0c, 32'hd7e13eaf, 1'h0)
`STIMULI(5'h0f, 5'h1c, 5'h0d, 32'h24343548, 1'h1)
`STIMULI(5'h1f, 5'h1c, 5'h0e, 32'hc645848c, 1'h1)
`STIMULI(5'h06, 5'h10, 5'h0f, 32'he2f310c5, 1'h1)
`STIMULI(5'h1a, 5'h00, 5'h10, 32'h39133172, 1'h1)
`STIMULI(5'h1e, 5'h15, 5'h11, 32'h28fc2151, 1'h1)
`STIMULI(5'h16, 5'h0a, 5'h12, 32'h3a9faf75, 1'h0)
`STIMULI(5'h13, 5'h1a, 5'h13, 32'h5ef0d9bd, 1'h1)
`STIMULI(5'h17, 5'h12, 5'h14, 32'hc9cec293, 1'h1)
`STIMULI(5'h13, 5'h0a, 5'h15, 32'h9639382c, 1'h1)
`STIMULI(5'h06, 5'h08, 5'h16, 32'h9a9aac35, 1'h0)
`STIMULI(5'h0b, 5'h15, 5'h17, 32'hc8a66691, 1'h1)
`STIMULI(5'h1a, 5'h0a, 5'h18, 32'h1e43493c, 1'h0)
`STIMULI(5'h1c, 5'h16, 5'h19, 32'h7b085df6, 1'h1)
`STIMULI(5'h1b, 5'h00, 5'h1a, 32'hc8ac2e91, 1'h1)
`STIMULI(5'h1c, 5'h18, 5'h1b, 32'h24de7d49, 1'h0)
`STIMULI(5'h03, 5'h12, 5'h1c, 32'h3631d56c, 1'h1)
`STIMULI(5'h1d, 5'h1f, 5'h1d, 32'h900b3620, 1'h0)
`STIMULI(5'h16, 5'h16, 5'h1e, 32'hc4fdac89, 1'h0)
`STIMULI(5'h1f, 5'h0f, 5'h1f, 32'h1e32a13c, 1'h0)
`STIMULI(5'h18, 5'h12, 5'h00, 32'hd6a13ead, 1'h0)
`STIMULI(5'h04, 5'h04, 5'h01, 32'hb62c246c, 1'h1)
`STIMULI(5'h13, 5'h19, 5'h02, 32'h32805765, 1'h0)
`STIMULI(5'h0a, 5'h16, 5'h03, 32'hbaaf1475, 1'h1)
`STIMULI(5'h1a, 5'h0f, 5'h04, 32'h575217ae, 1'h0)
`STIMULI(5'h14, 5'h02, 5'h05, 32'h04224f08, 1'h1)
`STIMULI(5'h0d, 5'h06, 5'h06, 32'he1c122c3, 1'h1)
`STIMULI(5'h05, 5'h0d, 5'h07, 32'h1a36dd34, 1'h0)
`STIMULI(5'h04, 5'h02, 5'h08, 32'hf7f2b4ef, 1'h0)
`STIMULI(5'h1a, 5'h17, 5'h09, 32'h06b5970d, 1'h1)
`STIMULI(5'h1a, 5'h13, 5'h0a, 32'hd57cc4aa, 1'h0)
`STIMULI(5'h09, 5'h14, 5'h0b, 32'hc1a7be83, 1'h1)
`STIMULI(5'h17, 5'h1d, 5'h0c, 32'h91132822, 1'h1)
`STIMULI(5'h13, 5'h12, 5'h0d, 32'h97c2a22f, 1'h1)
`STIMULI(5'h0a, 5'h1e, 5'h0e, 32'hf4f3b0e9, 1'h1)
`STIMULI(5'h14, 5'h0a, 5'h0f, 32'hb6be3c6d, 1'h0)
`STIMULI(5'h01, 5'h10, 5'h10, 32'h34d94969, 1'h1)
`STIMULI(5'h04, 5'h17, 5'h11, 32'h6ffed5df, 1'h1)
`STIMULI(5'h1a, 5'h0a, 5'h12, 32'h5ffe19bf, 1'h0)
`STIMULI(5'h16, 5'h15, 5'h13, 32'h70b99de1, 1'h1)
`STIMULI(5'h0d, 5'h06, 5'h14, 32'h1374a726, 1'h0)
`STIMULI(5'h1c, 5'h12, 5'h15, 32'h577c51ae, 1'h1)
`STIMULI(5'h1a, 5'h16, 5'h16, 32'h18dff531, 1'h1)
`STIMULI(5'h05, 5'h10, 5'h17, 32'h61bfdfc3, 1'h0)
`STIMULI(5'h10, 5'h1f, 5'h18, 32'hb7529a6e, 1'h1)
`STIMULI(5'h0e, 5'h1e, 5'h19, 32'h98edfc31, 1'h1)
`STIMULI(5'h0f, 5'h12, 5'h1a, 32'h77dcf5ef, 1'h0)
`STIMULI(5'h17, 5'h16, 5'h1b, 32'h9d01cc3a, 1'h0)
`STIMULI(5'h11, 5'h0d, 5'h1c, 32'h6d1237da, 1'h1)
`STIMULI(5'h0d, 5'h1e, 5'h1d, 32'h1bab7b37, 1'h0)
`STIMULI(5'h1b, 5'h1a, 5'h1e, 32'h9c8c8e39, 1'h0)
`STIMULI(5'h19, 5'h04, 5'h1f, 32'hdd9ee4bb, 1'h0)
`STIMULI(5'h06, 5'h1a, 5'h00, 32'h6b384dd6, 1'h0)
`STIMULI(5'h0e, 5'h1c, 5'h01, 32'h48753190, 1'h1)
`STIMULI(5'h14, 5'h07, 5'h02, 32'hd0edf8a1, 1'h1)
`STIMULI(5'h18, 5'h07, 5'h03, 32'hf2496ee4, 1'h1)
`STIMULI(5'h15, 5'h04, 5'h04, 32'h0da3751b, 1'h0)
`STIMULI(5'h17, 5'h17, 5'h05, 32'h9cf84039, 1'h0)
`STIMULI(5'h10, 5'h0f, 5'h06, 32'h923c2224, 1'h1)
`STIMULI(5'h11, 5'h0f, 5'h07, 32'h51aa6da3, 1'h0)
`STIMULI(5'h1c, 5'h13, 5'h08, 32'h38bfff71, 1'h0)
`STIMULI(5'h0d, 5'h15, 5'h09, 32'h92128e24, 1'h0)
`STIMULI(5'h0b, 5'h08, 5'h0a, 32'hb381c267, 1'h1)
`STIMULI(5'h0c, 5'h03, 5'h0b, 32'h5b85a5b7, 1'h0)
`STIMULI(5'h0c, 5'h13, 5'h0c, 32'hb87c0070, 1'h0)
`STIMULI(5'h12, 5'h1c, 5'h0d, 32'h38d6bf71, 1'h1)
`STIMULI(5'h1a, 5'h17, 5'h0e, 32'hcded4a9b, 1'h0)
`STIMULI(5'h10, 5'h07, 5'h0f, 32'h8a9d9815, 1'h0)
`STIMULI(5'h1e, 5'h1b, 5'h10, 32'h2efb4f5d, 1'h0)
`STIMULI(5'h05, 5'h02, 5'h11, 32'hb2503664, 1'h1)
`STIMULI(5'h05, 5'h06, 5'h12, 32'hf2e4f2e5, 1'h0)
`STIMULI(5'h06, 5'h0d, 5'h13, 32'h9b578e36, 1'h1)
`STIMULI(5'h08, 5'h06, 5'h14, 32'he70b7cce, 1'h1)
`STIMULI(5'h11, 5'h12, 5'h15, 32'h66071bcc, 1'h1)
`STIMULI(5'h15, 5'h1a, 5'h16, 32'h53daada7, 1'h1)
`STIMULI(5'h0f, 5'h16, 5'h17, 32'h6b1f87d6, 1'h0)
`STIMULI(5'h1d, 5'h06, 5'h18, 32'h9e57de3c, 1'h0)
`STIMULI(5'h0f, 5'h14, 5'h19, 32'h9b444c36, 1'h1)
`STIMULI(5'h0b, 5'h1e, 5'h1a, 32'h53e02ba7, 1'h1)
`STIMULI(5'h18, 5'h02, 5'h1b, 32'h148c4b29, 1'h0)
`STIMULI(5'h1d, 5'h1e, 5'h1c, 32'h1b5d8736, 1'h1)
`STIMULI(5'h16, 5'h1e, 5'h1d, 32'hd91570b2, 1'h0)
`STIMULI(5'h0b, 5'h04, 5'h1e, 32'h36fae36d, 1'h0)
`STIMULI(5'h09, 5'h06, 5'h1f, 32'h8c435818, 1'h1)
`STIMULI(5'h02, 5'h03, 5'h00, 32'h231f4d46, 1'h0)
`STIMULI(5'h1f, 5'h14, 5'h01, 32'h3110eb62, 1'h1)
`STIMULI(5'h08, 5'h09, 5'h02, 32'h633809c6, 1'h1)
`STIMULI(5'h0e, 5'h1b, 5'h03, 32'hc29cf885, 1'h1)
`STIMULI(5'h05, 5'h18, 5'h04, 32'h2299c145, 1'h1)
`STIMULI(5'h0b, 5'h0c, 5'h05, 32'h58d9e1b1, 1'h1)
`STIMULI(5'h12, 5'h14, 5'h06, 32'he78090cf, 1'h1)
`STIMULI(5'h05, 5'h08, 5'h07, 32'h0e082d1c, 1'h0)
`STIMULI(5'h1c, 5'h1a, 5'h08, 32'h9ff7383f, 1'h1)
`STIMULI(5'h11, 5'h03, 5'h09, 32'h3664356c, 1'h0)
`STIMULI(5'h12, 5'h16, 5'h0a, 32'hbc2d2e78, 1'h1)
`STIMULI(5'h10, 5'h1c, 5'h0b, 32'h622ebbc4, 1'h0)
`STIMULI(5'h1a, 5'h1e, 5'h0c, 32'h4783c98f, 1'h1)
`STIMULI(5'h16, 5'h0a, 5'h0d, 32'h42f88d85, 1'h0)
`STIMULI(5'h01, 5'h15, 5'h0e, 32'hf15a56e2, 1'h1)
`STIMULI(5'h06, 5'h1f, 5'h0f, 32'h97d9242f, 1'h1)
`STIMULI(5'h13, 5'h0b, 5'h10, 32'h28614550, 1'h1)
`STIMULI(5'h06, 5'h1b, 5'h11, 32'he8f84ad1, 1'h0)
`STIMULI(5'h13, 5'h1c, 5'h12, 32'hbefc3c7d, 1'h1)
`STIMULI(5'h17, 5'h15, 5'h13, 32'hc992b093, 1'h0)
`STIMULI(5'h1d, 5'h14, 5'h14, 32'h74fb41e9, 1'h1)
`STIMULI(5'h08, 5'h11, 5'h15, 32'hc0619280, 1'h0)
`STIMULI(5'h0f, 5'h0d, 5'h16, 32'h2ab2d355, 1'h0)
`STIMULI(5'h16, 5'h05, 5'h17, 32'h890d5e12, 1'h0)
`STIMULI(5'h19, 5'h08, 5'h18, 32'hdb3b10b6, 1'h1)
`STIMULI(5'h12, 5'h14, 5'h19, 32'h4e134b9c, 1'h1)
`STIMULI(5'h10, 5'h0f, 5'h1a, 32'hb75dd06e, 1'h1)
`STIMULI(5'h11, 5'h18, 5'h1b, 32'h7145f9e2, 1'h0)
`STIMULI(5'h14, 5'h03, 5'h1c, 32'h487bc790, 1'h1)
`STIMULI(5'h1b, 5'h1c, 5'h1d, 32'ha9d11453, 1'h0)
`STIMULI(5'h03, 5'h1f, 5'h1e, 32'h5270a7a4, 1'h0)
`STIMULI(5'h16, 5'h19, 5'h1f, 32'h5967fdb2, 1'h1)
`STIMULI(5'h19, 5'h13, 5'h00, 32'had3e3a5a, 1'h1)
`STIMULI(5'h19, 5'h1e, 5'h01, 32'h2f07575e, 1'h0)
`STIMULI(5'h15, 5'h17, 5'h02, 32'h73068be6, 1'h0)
`STIMULI(5'h1c, 5'h12, 5'h03, 32'h2c71b358, 1'h1)
`STIMULI(5'h0c, 5'h06, 5'h04, 32'h149cfd29, 1'h0)
`STIMULI(5'h02, 5'h14, 5'h05, 32'h1c4f3338, 1'h1)
`STIMULI(5'h16, 5'h0b, 5'h06, 32'h1eb6713d, 1'h0)
`STIMULI(5'h08, 5'h04, 5'h07, 32'h29981d53, 1'h0)
`STIMULI(5'h09, 5'h1e, 5'h08, 32'h23806347, 1'h1)
`STIMULI(5'h17, 5'h08, 5'h09, 32'hc5b28c8b, 1'h1)
`STIMULI(5'h1c, 5'h02, 5'h0a, 32'h48270d90, 1'h1)
`STIMULI(5'h01, 5'h04, 5'h0b, 32'h116b0122, 1'h1)
`STIMULI(5'h1a, 5'h1b, 5'h0c, 32'hd39282a7, 1'h1)
`STIMULI(5'h1c, 5'h06, 5'h0d, 32'hbdb00a7b, 1'h0)
`STIMULI(5'h07, 5'h1b, 5'h0e, 32'hbb62d276, 1'h1)
`STIMULI(5'h1b, 5'h04, 5'h0f, 32'h83b8e007, 1'h0)
`STIMULI(5'h1d, 5'h02, 5'h10, 32'hfdf32cfb, 1'h0)
`STIMULI(5'h07, 5'h1f, 5'h11, 32'h18ff0f31, 1'h1)
`STIMULI(5'h17, 5'h1e, 5'h12, 32'h8bebf617, 1'h0)
`STIMULI(5'h14, 5'h1a, 5'h13, 32'h92330224, 1'h0)
`STIMULI(5'h1b, 5'h09, 5'h14, 32'h09abf513, 1'h1)
`STIMULI(5'h10, 5'h0e, 5'h15, 32'hb113bc62, 1'h1)
`STIMULI(5'h14, 5'h04, 5'h16, 32'hb8906a71, 1'h0)
`STIMULI(5'h1d, 5'h15, 5'h17, 32'h4bd16997, 1'h0)
`STIMULI(5'h17, 5'h04, 5'h18, 32'hd1e432a3, 1'h0)
`STIMULI(5'h06, 5'h0f, 5'h19, 32'h0962fb12, 1'h1)
`STIMULI(5'h18, 5'h06, 5'h1a, 32'h78fde7f1, 1'h0)
`STIMULI(5'h0d, 5'h0a, 5'h1b, 32'hc4f6d689, 1'h1)
`STIMULI(5'h19, 5'h14, 5'h1c, 32'h97d4f82f, 1'h1)
`STIMULI(5'h19, 5'h0e, 5'h1d, 32'h3b666b76, 1'h0)
`STIMULI(5'h16, 5'h09, 5'h1e, 32'h6915dbd2, 1'h1)
`STIMULI(5'h04, 5'h1a, 5'h1f, 32'he054d0c0, 1'h1)
`STIMULI(5'h13, 5'h08, 5'h00, 32'h947d1828, 1'h0)
`STIMULI(5'h17, 5'h01, 5'h01, 32'h0d60711a, 1'h1)
`STIMULI(5'h1b, 5'h00, 5'h02, 32'h86017c0c, 1'h1)
`STIMULI(5'h0a, 5'h06, 5'h03, 32'hdc8f9cb9, 1'h1)
`STIMULI(5'h04, 5'h06, 5'h04, 32'h7e152bfc, 1'h0)
`STIMULI(5'h04, 5'h1c, 5'h05, 32'h17e0332f, 1'h0)
`STIMULI(5'h16, 5'h04, 5'h06, 32'hb105c062, 1'h1)
`STIMULI(5'h1a, 5'h05, 5'h07, 32'h6aa23fd5, 1'h1)
`STIMULI(5'h01, 5'h19, 5'h08, 32'h15437f2a, 1'h0)
`STIMULI(5'h09, 5'h03, 5'h09, 32'h9e05923c, 1'h1)
`STIMULI(5'h0e, 5'h0b, 5'h0a, 32'h2c175b58, 1'h0)
`STIMULI(5'h08, 5'h19, 5'h0b, 32'hd10276a2, 1'h1)
`STIMULI(5'h1b, 5'h1d, 5'h0c, 32'h8e102a1c, 1'h1)
`STIMULI(5'h1f, 5'h12, 5'h0d, 32'h7c8537f9, 1'h1)
`STIMULI(5'h0b, 5'h08, 5'h0e, 32'h442ebf88, 1'h1)
`STIMULI(5'h0e, 5'h1f, 5'h0f, 32'h5f84cdbf, 1'h0)
`STIMULI(5'h10, 5'h1b, 5'h10, 32'h689903d1, 1'h0)
`STIMULI(5'h1f, 5'h03, 5'h11, 32'h536c81a6, 1'h0)
`STIMULI(5'h1c, 5'h18, 5'h12, 32'h1d5c1f3a, 1'h1)
`STIMULI(5'h03, 5'h00, 5'h13, 32'h38008570, 1'h1)
`STIMULI(5'h0a, 5'h17, 5'h14, 32'h0d859b1b, 1'h1)
`STIMULI(5'h0e, 5'h01, 5'h15, 32'hcea5949d, 1'h1)
`STIMULI(5'h0c, 5'h09, 5'h16, 32'h549b73a9, 1'h1)
`STIMULI(5'h00, 5'h16, 5'h17, 32'h2fb3a15f, 1'h0)
`STIMULI(5'h1f, 5'h13, 5'h18, 32'h423b4584, 1'h0)
`STIMULI(5'h0e, 5'h10, 5'h19, 32'hb13b5862, 1'h0)
`STIMULI(5'h13, 5'h1d, 5'h1a, 32'heb686ad6, 1'h0)
`STIMULI(5'h0e, 5'h01, 5'h1b, 32'h4d66e59a, 1'h1)
`STIMULI(5'h09, 5'h01, 5'h1c, 32'h48d11991, 1'h0)
`STIMULI(5'h04, 5'h02, 5'h1d, 32'h075d6f0e, 1'h0)
`STIMULI(5'h10, 5'h1d, 5'h1e, 32'hb1127e62, 1'h1)
`STIMULI(5'h09, 5'h1f, 5'h1f, 32'h2851d550, 1'h0)
`STIMULI(5'h11, 5'h19, 5'h00, 32'h3fc3e97f, 1'h0)
`STIMULI(5'h0b, 5'h1f, 5'h01, 32'ha3243c46, 1'h1)
`STIMULI(5'h10, 5'h0c, 5'h02, 32'h1dd0df3b, 1'h1)
`STIMULI(5'h18, 5'h05, 5'h03, 32'h2bbeb757, 1'h0)
`STIMULI(5'h00, 5'h04, 5'h04, 32'h156a472a, 1'h1)
`STIMULI(5'h15, 5'h06, 5'h05, 32'hc814e490, 1'h0)
`STIMULI(5'h05, 5'h05, 5'h06, 32'h539681a7, 1'h1)
`STIMULI(5'h11, 5'h06, 5'h07, 32'h836e8e06, 1'h0)
`STIMULI(5'h1b, 5'h00, 5'h08, 32'h23288946, 1'h1)
`STIMULI(5'h07, 5'h0b, 5'h09, 32'ha9654a52, 1'h0)
`STIMULI(5'h05, 5'h05, 5'h0a, 32'hb8a61871, 1'h0)
`STIMULI(5'h02, 5'h12, 5'h0b, 32'h34bd1d69, 1'h0)
`STIMULI(5'h07, 5'h0e, 5'h0c, 32'h4464c388, 1'h0)
`STIMULI(5'h0c, 5'h07, 5'h0d, 32'h1f00153e, 1'h0)
`STIMULI(5'h05, 5'h0f, 5'h0e, 32'h5fe61bbf, 1'h0)
`STIMULI(5'h13, 5'h11, 5'h0f, 32'ha884e851, 1'h1)
`STIMULI(5'h17, 5'h08, 5'h10, 32'hfd3ac8fa, 1'h0)
`STIMULI(5'h1b, 5'h12, 5'h11, 32'hb548a46a, 1'h1)
`STIMULI(5'h05, 5'h0f, 5'h12, 32'h32f4b965, 1'h0)
`STIMULI(5'h1f, 5'h03, 5'h13, 32'ha9c33653, 1'h0)
`STIMULI(5'h07, 5'h06, 5'h14, 32'h04f02f09, 1'h1)
`STIMULI(5'h1f, 5'h19, 5'h15, 32'hfb9f1ef7, 1'h0)
`STIMULI(5'h14, 5'h1e, 5'h16, 32'h91fbea23, 1'h0)
`STIMULI(5'h10, 5'h0d, 5'h17, 32'h9cfc0839, 1'h1)
`STIMULI(5'h14, 5'h05, 5'h18, 32'h48284990, 1'h1)
`STIMULI(5'h08, 5'h19, 5'h19, 32'hb5a4686b, 1'h0)
`STIMULI(5'h0b, 5'h07, 5'h1a, 32'hdd4560ba, 1'h0)
`STIMULI(5'h0f, 5'h1f, 5'h1b, 32'h745e23e8, 1'h1)
`STIMULI(5'h19, 5'h11, 5'h1c, 32'h36d8296d, 1'h0)
`STIMULI(5'h06, 5'h1d, 5'h1d, 32'h533e25a6, 1'h0)
`STIMULI(5'h16, 5'h0b, 5'h1e, 32'h1c8e9339, 1'h0)
`STIMULI(5'h19, 5'h14, 5'h1f, 32'ha4a70849, 1'h1)
`STIMULI(5'h09, 5'h15, 5'h00, 32'hf1faa6e3, 1'h0)
`STIMULI(5'h01, 5'h10, 5'h01, 32'hd35ab6a6, 1'h0)
`STIMULI(5'h04, 5'h1c, 5'h02, 32'hb81cb070, 1'h0)
`STIMULI(5'h00, 5'h18, 5'h03, 32'h1ec7013d, 1'h0)
`STIMULI(5'h0b, 5'h05, 5'h04, 32'had04525a, 1'h0)
`STIMULI(5'h0e, 5'h0e, 5'h05, 32'hf57544ea, 1'h1)
`STIMULI(5'h0c, 5'h0d, 5'h06, 32'hf790b0ef, 1'h1)
`STIMULI(5'h1e, 5'h1b, 5'h07, 32'h12450f24, 1'h0)
`STIMULI(5'h02, 5'h1f, 5'h08, 32'h571783ae, 1'h1)
`STIMULI(5'h0a, 5'h0d, 5'h09, 32'h5dd9b3bb, 1'h1)
`STIMULI(5'h16, 5'h00, 5'h0a, 32'hba7b4674, 1'h0)
`STIMULI(5'h06, 5'h1d, 5'h0b, 32'hfc62f2f8, 1'h0)
`STIMULI(5'h1f, 5'h14, 5'h0c, 32'h5ff84dbf, 1'h0)
`STIMULI(5'h0d, 5'h17, 5'h0d, 32'h10a8a121, 1'h0)
`STIMULI(5'h06, 5'h1e, 5'h0e, 32'h9eb0e43d, 1'h0)
`STIMULI(5'h18, 5'h13, 5'h0f, 32'h48013590, 1'h0)
`STIMULI(5'h15, 5'h13, 5'h10, 32'h2cc08159, 1'h0)
`STIMULI(5'h03, 5'h11, 5'h11, 32'h679b77cf, 1'h1)
`STIMULI(5'h0e, 5'h1d, 5'h12, 32'h885dc210, 1'h1)
`STIMULI(5'h1d, 5'h16, 5'h13, 32'h82431804, 1'h0)
`STIMULI(5'h09, 5'h18, 5'h14, 32'h9053b220, 1'h0)
`STIMULI(5'h1b, 5'h1f, 5'h15, 32'h668859cd, 1'h1)
`STIMULI(5'h02, 5'h1e, 5'h16, 32'h3fd9d37f, 1'h1)
`STIMULI(5'h1b, 5'h1a, 5'h17, 32'he7f2a0cf, 1'h1)
`STIMULI(5'h0f, 5'h03, 5'h18, 32'h5b933bb7, 1'h1)
`STIMULI(5'h09, 5'h06, 5'h19, 32'h12a62725, 1'h0)
`STIMULI(5'h01, 5'h0c, 5'h1a, 32'h993cc632, 1'h0)
`STIMULI(5'h01, 5'h1f, 5'h1b, 32'hcfa4909f, 1'h0)
`STIMULI(5'h16, 5'h02, 5'h1c, 32'hd9522ab2, 1'h0)
`STIMULI(5'h05, 5'h1d, 5'h1d, 32'h30908b61, 1'h1)
`STIMULI(5'h04, 5'h1b, 5'h1e, 32'h59b215b3, 1'h0)
`STIMULI(5'h1d, 5'h1f, 5'h1f, 32'h349c6d69, 1'h1)
`STIMULI(5'h0c, 5'h00, 5'h00, 32'hca095494, 1'h0)
`STIMULI(5'h1b, 5'h05, 5'h01, 32'h8d0be21a, 1'h1)
`STIMULI(5'h1e, 5'h06, 5'h02, 32'hce8cf09d, 1'h1)
`STIMULI(5'h10, 5'h1f, 5'h03, 32'h66707bcc, 1'h1)
`STIMULI(5'h08, 5'h06, 5'h04, 32'h334b5166, 1'h1)
`STIMULI(5'h00, 5'h09, 5'h05, 32'hb4895669, 1'h1)
`STIMULI(5'h0d, 5'h13, 5'h06, 32'hca1c5094, 1'h0)
`STIMULI(5'h07, 5'h0e, 5'h07, 32'ha16dbe42, 1'h1)
`STIMULI(5'h1d, 5'h1c, 5'h08, 32'h16f86f2d, 1'h0)
`STIMULI(5'h03, 5'h11, 5'h09, 32'hbd6ac87a, 1'h1)
`STIMULI(5'h0f, 5'h00, 5'h0a, 32'h7a3ee3f4, 1'h1)
`STIMULI(5'h01, 5'h1f, 5'h0b, 32'h13bbf927, 1'h1)
`STIMULI(5'h1a, 5'h08, 5'h0c, 32'he632c4cc, 1'h0)
`STIMULI(5'h00, 5'h0b, 5'h0d, 32'h8906de12, 1'h0)
`STIMULI(5'h15, 5'h19, 5'h0e, 32'h4cb72199, 1'h1)
`STIMULI(5'h03, 5'h16, 5'h0f, 32'h9341b026, 1'h1)
`STIMULI(5'h06, 5'h1f, 5'h10, 32'h44122788, 1'h0)
`STIMULI(5'h16, 5'h1d, 5'h11, 32'h9f6cfa3e, 1'h1)
`STIMULI(5'h08, 5'h17, 5'h12, 32'hd53f3caa, 1'h1)
`STIMULI(5'h09, 5'h06, 5'h13, 32'h08482b10, 1'h0)
`STIMULI(5'h1f, 5'h06, 5'h14, 32'h6c1829d8, 1'h0)
`STIMULI(5'h0e, 5'h10, 5'h15, 32'h89e94013, 1'h1)
`STIMULI(5'h04, 5'h1d, 5'h16, 32'h695d29d2, 1'h1)
`STIMULI(5'h03, 5'h14, 5'h17, 32'h50df69a1, 1'h0)
`STIMULI(5'h02, 5'h0d, 5'h18, 32'h50641da0, 1'h0)
`STIMULI(5'h1d, 5'h09, 5'h19, 32'h504897a0, 1'h1)
`STIMULI(5'h0e, 5'h0e, 5'h1a, 32'he5f69ccb, 1'h0)
`STIMULI(5'h0f, 5'h13, 5'h1b, 32'h21022f42, 1'h1)
`STIMULI(5'h04, 5'h0d, 5'h1c, 32'h43a71b87, 1'h0)
`STIMULI(5'h1b, 5'h16, 5'h1d, 32'h7cdc9ff9, 1'h1)
`STIMULI(5'h0d, 5'h10, 5'h1e, 32'hd2a508a5, 1'h1)
`STIMULI(5'h15, 5'h1d, 5'h1f, 32'h237a0346, 1'h0)
`STIMULI(5'h00, 5'h1b, 5'h00, 32'hc2d7f285, 1'h1)
`STIMULI(5'h15, 5'h05, 5'h01, 32'hcb3fbe96, 1'h1)
`STIMULI(5'h1c, 5'h1b, 5'h02, 32'hd6c9a2ad, 1'h1)
`STIMULI(5'h11, 5'h12, 5'h03, 32'h5f8325bf, 1'h1)
`STIMULI(5'h11, 5'h1e, 5'h04, 32'hb2a73c65, 1'h1)
`STIMULI(5'h15, 5'h00, 5'h05, 32'h65d917cb, 1'h1)
`STIMULI(5'h02, 5'h05, 5'h06, 32'h34615f68, 1'h1)
`STIMULI(5'h0c, 5'h03, 5'h07, 32'ha7309e4e, 1'h0)
`STIMULI(5'h0a, 5'h11, 5'h08, 32'h24b34949, 1'h1)
`STIMULI(5'h1b, 5'h15, 5'h09, 32'h562091ac, 1'h1)
`STIMULI(5'h14, 5'h03, 5'h0a, 32'hbc98f079, 1'h1)
`STIMULI(5'h1b, 5'h17, 5'h0b, 32'h92902e25, 1'h1)
`STIMULI(5'h09, 5'h1e, 5'h0c, 32'h787c2df0, 1'h1)
`STIMULI(5'h1e, 5'h06, 5'h0d, 32'h8ba2ca17, 1'h0)
`STIMULI(5'h13, 5'h1d, 5'h0e, 32'h7220cde4, 1'h1)
`STIMULI(5'h0f, 5'h03, 5'h0f, 32'h4b8e5f97, 1'h1)
`STIMULI(5'h1d, 5'h06, 5'h10, 32'h6c17bdd8, 1'h1)
`STIMULI(5'h0b, 5'h0a, 5'h11, 32'h9dc52c3b, 1'h1)
`STIMULI(5'h00, 5'h09, 5'h12, 32'hcd41269a, 1'h0)
`STIMULI(5'h08, 5'h18, 5'h13, 32'h2e9a6d5d, 1'h0)
`STIMULI(5'h0f, 5'h02, 5'h14, 32'h70a58de1, 1'h1)
`STIMULI(5'h1f, 5'h07, 5'h15, 32'h2c49db58, 1'h1)
`STIMULI(5'h01, 5'h05, 5'h16, 32'h55adf1ab, 1'h0)
`STIMULI(5'h03, 5'h0b, 5'h17, 32'h040a6108, 1'h1)
`STIMULI(5'h16, 5'h1b, 5'h18, 32'h5682f1ad, 1'h1)
`STIMULI(5'h08, 5'h0b, 5'h19, 32'h8293b405, 1'h0)
`STIMULI(5'h02, 5'h08, 5'h1a, 32'h061ae30c, 1'h1)
`STIMULI(5'h1c, 5'h05, 5'h1b, 32'h563efdac, 1'h0)
`STIMULI(5'h1f, 5'h01, 5'h1c, 32'h253efb4a, 1'h1)
`STIMULI(5'h1d, 5'h18, 5'h1d, 32'he1aa64c3, 1'h0)
`STIMULI(5'h1e, 5'h01, 5'h1e, 32'had8f6c5b, 1'h1)
`STIMULI(5'h1b, 5'h02, 5'h1f, 32'h2887c751, 1'h0)
`STIMULI(5'h05, 5'h1a, 5'h00, 32'hb34e8266, 1'h0)
`STIMULI(5'h01, 5'h13, 5'h01, 32'h94fe4829, 1'h0)
`STIMULI(5'h16, 5'h03, 5'h02, 32'h427ac584, 1'h0)
`STIMULI(5'h04, 5'h00, 5'h03, 32'h12c70125, 1'h0)
`STIMULI(5'h18, 5'h19, 5'h04, 32'h518019a3, 1'h0)
`STIMULI(5'h10, 5'h19, 5'h05, 32'hb5ec886b, 1'h0)
`STIMULI(5'h1e, 5'h0b, 5'h06, 32'hdb87deb7, 1'h0)
`STIMULI(5'h05, 5'h15, 5'h07, 32'h85d5ae0b, 1'h1)
`STIMULI(5'h1e, 5'h14, 5'h08, 32'h9e30123c, 1'h1)
`STIMULI(5'h12, 5'h0f, 5'h09, 32'h42030784, 1'h0)
`STIMULI(5'h02, 5'h00, 5'h0a, 32'hc2316e84, 1'h1)
`STIMULI(5'h11, 5'h1a, 5'h0b, 32'hbca79679, 1'h0)
`STIMULI(5'h16, 5'h01, 5'h0c, 32'h543c85a8, 1'h0)
`STIMULI(5'h17, 5'h00, 5'h0d, 32'he80468d0, 1'h1)
`STIMULI(5'h17, 5'h1f, 5'h0e, 32'hd315e8a6, 1'h1)
`STIMULI(5'h13, 5'h1c, 5'h0f, 32'h9e2f3a3c, 1'h1)
`STIMULI(5'h07, 5'h1a, 5'h10, 32'ha9b94253, 1'h1)
`STIMULI(5'h10, 5'h05, 5'h11, 32'hafac105f, 1'h0)
`STIMULI(5'h19, 5'h17, 5'h12, 32'h200b8140, 1'h0)
`STIMULI(5'h15, 5'h06, 5'h13, 32'h9401de28, 1'h0)
`STIMULI(5'h17, 5'h15, 5'h14, 32'h9263e024, 1'h1)
`STIMULI(5'h0a, 5'h10, 5'h15, 32'h603223c0, 1'h1)
`STIMULI(5'h17, 5'h19, 5'h16, 32'h87f4280f, 1'h1)
`STIMULI(5'h0f, 5'h05, 5'h17, 32'h19bb8933, 1'h0)
`STIMULI(5'h0d, 5'h1d, 5'h18, 32'hf9d7b2f3, 1'h0)
`STIMULI(5'h09, 5'h11, 5'h19, 32'h498f8593, 1'h0)
`STIMULI(5'h07, 5'h0b, 5'h1a, 32'hb8519670, 1'h1)
`STIMULI(5'h01, 5'h16, 5'h1b, 32'h8922fa12, 1'h0)
`STIMULI(5'h1c, 5'h05, 5'h1c, 32'hc981cc93, 1'h1)
`STIMULI(5'h16, 5'h07, 5'h1d, 32'hd481d8a9, 1'h0)
`STIMULI(5'h1a, 5'h1f, 5'h1e, 32'hcc994099, 1'h1)
`STIMULI(5'h01, 5'h1c, 5'h1f, 32'h670dbbce, 1'h1)
`STIMULI(5'h14, 5'h0d, 5'h00, 32'h4e55019c, 1'h0)
`STIMULI(5'h09, 5'h05, 5'h01, 32'hfd4f84fa, 1'h1)
`STIMULI(5'h1c, 5'h1d, 5'h02, 32'h7f4857fe, 1'h1)
`STIMULI(5'h01, 5'h13, 5'h03, 32'h35040b6a, 1'h0)
`STIMULI(5'h08, 5'h1c, 5'h04, 32'h523de5a4, 1'h1)
`STIMULI(5'h0a, 5'h0e, 5'h05, 32'h9d4baa3a, 1'h1)
`STIMULI(5'h0a, 5'h03, 5'h06, 32'ha0b7ce41, 1'h0)
`STIMULI(5'h1f, 5'h16, 5'h07, 32'h8ba4ee17, 1'h0)
`STIMULI(5'h06, 5'h10, 5'h08, 32'hfd56cefa, 1'h0)
`STIMULI(5'h01, 5'h0f, 5'h09, 32'h271a2f4e, 1'h0)
`STIMULI(5'h0f, 5'h04, 5'h0a, 32'h47b05d8f, 1'h1)
`STIMULI(5'h1a, 5'h18, 5'h0b, 32'h01ca2d03, 1'h0)
`STIMULI(5'h1f, 5'h15, 5'h0c, 32'h52dbcfa5, 1'h0)
`STIMULI(5'h11, 5'h0b, 5'h0d, 32'h39b3b573, 1'h0)
`STIMULI(5'h13, 5'h0c, 5'h0e, 32'hefbe74df, 1'h0)
`STIMULI(5'h1d, 5'h18, 5'h0f, 32'h246c4748, 1'h0)
`STIMULI(5'h06, 5'h05, 5'h10, 32'hdddebabb, 1'h0)
`STIMULI(5'h0d, 5'h13, 5'h11, 32'h2e29a35c, 1'h0)
`STIMULI(5'h0d, 5'h1c, 5'h12, 32'h794649f2, 1'h1)
`STIMULI(5'h06, 5'h05, 5'h13, 32'h83468006, 1'h1)
`STIMULI(5'h0f, 5'h01, 5'h14, 32'he1bb26c3, 1'h1)
`STIMULI(5'h07, 5'h16, 5'h15, 32'h842a1c08, 1'h0)
`STIMULI(5'h1b, 5'h13, 5'h16, 32'hbf57d07e, 1'h1)
`STIMULI(5'h12, 5'h01, 5'h17, 32'h963ae02c, 1'h1)
`STIMULI(5'h00, 5'h1d, 5'h18, 32'h224a6544, 1'h0)
`STIMULI(5'h13, 5'h14, 5'h19, 32'hd14404a2, 1'h0)
`STIMULI(5'h1f, 5'h01, 5'h1a, 32'h3742bd6e, 1'h1)
`STIMULI(5'h11, 5'h01, 5'h1b, 32'hff7628fe, 1'h0)
`STIMULI(5'h09, 5'h18, 5'h1c, 32'h17d78d2f, 1'h0)
`STIMULI(5'h0b, 5'h01, 5'h1d, 32'h96eafe2d, 1'h0)
`STIMULI(5'h1f, 5'h13, 5'h1e, 32'hcdea849b, 1'h0)
`STIMULI(5'h0f, 5'h10, 5'h1f, 32'h6e53dfdc, 1'h0)
`STIMULI(5'h1b, 5'h1a, 5'h00, 32'h22d36f45, 1'h1)
`STIMULI(5'h11, 5'h0e, 5'h01, 32'h233b6f46, 1'h0)
`STIMULI(5'h13, 5'h02, 5'h02, 32'hf6da58ed, 1'h0)
`STIMULI(5'h18, 5'h0a, 5'h03, 32'h2702454e, 1'h0)
`STIMULI(5'h03, 5'h06, 5'h04, 32'h1348a326, 1'h1)
`STIMULI(5'h15, 5'h13, 5'h05, 32'h607e7bc0, 1'h1)
`STIMULI(5'h09, 5'h05, 5'h06, 32'ha1192e42, 1'h1)
`STIMULI(5'h04, 5'h13, 5'h07, 32'hf2e65ee5, 1'h1)
`STIMULI(5'h08, 5'h0b, 5'h08, 32'h180f7930, 1'h1)
`STIMULI(5'h1a, 5'h1a, 5'h09, 32'h376e056e, 1'h1)
`STIMULI(5'h07, 5'h14, 5'h0a, 32'h85bdba0b, 1'h1)
`STIMULI(5'h04, 5'h15, 5'h0b, 32'hfdbff2fb, 1'h1)
`STIMULI(5'h1f, 5'h15, 5'h0c, 32'he9c206d3, 1'h1)
`STIMULI(5'h0e, 5'h11, 5'h0d, 32'he838b2d0, 1'h0)
`STIMULI(5'h0d, 5'h08, 5'h0e, 32'h04426f08, 1'h1)
`STIMULI(5'h10, 5'h0b, 5'h0f, 32'he38d82c7, 1'h0)
`STIMULI(5'h17, 5'h0a, 5'h10, 32'hc570208a, 1'h0)
`STIMULI(5'h1f, 5'h10, 5'h11, 32'h7e45e7fc, 1'h1)
`STIMULI(5'h0f, 5'h0b, 5'h12, 32'h80998201, 1'h1)
`STIMULI(5'h06, 5'h02, 5'h13, 32'hf33052e6, 1'h1)
`STIMULI(5'h05, 5'h1d, 5'h14, 32'h8b135a16, 1'h0)
`STIMULI(5'h03, 5'h15, 5'h15, 32'h42b9c585, 1'h0)
`STIMULI(5'h1b, 5'h07, 5'h16, 32'hf700e8ee, 1'h1)
`STIMULI(5'h10, 5'h16, 5'h17, 32'h69d069d3, 1'h0)
`STIMULI(5'h01, 5'h19, 5'h18, 32'h13c30927, 1'h0)
`STIMULI(5'h14, 5'h07, 5'h19, 32'hd1b932a3, 1'h1)
`STIMULI(5'h01, 5'h0b, 5'h1a, 32'h39965373, 1'h0)
`STIMULI(5'h17, 5'h18, 5'h1b, 32'h2b008756, 1'h0)
`STIMULI(5'h08, 5'h12, 5'h1c, 32'h93a83c27, 1'h0)
`STIMULI(5'h16, 5'h1b, 5'h1d, 32'h366dd36c, 1'h0)
`STIMULI(5'h1f, 5'h1f, 5'h1e, 32'h0bab3717, 1'h0)
